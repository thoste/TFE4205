��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8FΣ�?����ǝ��.�mF�q�TCђQ���hcX~�`&
?qA�$�#Vǜ��O��a�Fo[������2�do�\�IG4T��(��ٕ(J%��ͦ��b}�OI�Rg x�sL���,�yۨTD�wxN�1��ؿA�T��ǹ�=��[���N�n��s�:�E�6�e�0�b����嵱�Sݩ"��(�Q ����Ɣ��CS��Gn@1�F�i�X=Nn�$��a�߃����Z�C)�y��;u}S���Uһ���?1c��y��t�,���%nd���cj�\�����f��:��u��zg9o���b�>�̶�J�e��+��[�ƕ2���X�*팆��W�SW�ZiL�-�Dm� ��}'.c��v�t�τs�5X��V��	8�B� `4�oY��T$��-��n{j����9���Ior0���
L��1��8�6A5.+��0�,y$�&!a �_Z���n݆bb�����Q���`n=9�Rq���Gw�.%����>���J����P5��U�=��	\-�N�Ҁ�5����y޺$�(8�,���׵7;�/�W �wE�t�,n�ɘ�s�/em�>�H.��A�W��a�.�x�����Man�(�j�����r����&{,��^���C�z��Ht��wb悡l���{yۗ�v�����g��f�MW��΃�fy:�8Ny�1�.1<ۧ�#���Ð�����P��^�p/�������r|�E��!4�T�Js��u
:�s�7z�R؏��9\|�O��*QF��~
9���:�g�Ӎ�S]l��xC�`y��2׼�IQ���"�PX���ť��q��N'�Mh�k����)��?%e��4K5#qg�������إ�u�|O����������}�#�&l�e�z�n�64	�?�cCBٗf����I��W�n���0���Y��1�_*ƣ�V�w�z�2��@2)�����o�6���2fݲZ���4����s/ۭ?u3���AY�`�"ܕa��ӷ����W����gI���=T5e��� �*B�a���:����v��⸎�3���r�8{���)K'�s���FP�@�v�G[ȇ�-��7��7(~n�a(y,�+c�����icO�l�C�+=��N��H˾T%슗�"<7�#�^{�����e�7&.IP\+�ӈ}}��z��E&��^�WE��)ԔE`*�ZV}E(��95��<<#b�*�r$J�Bl��I�z���ڶ�HI�
�ڗW|�Z�J������*�I�~'�����v��:�Y~���m)�]{O����d\���+ �ɓo�ƀ�qc��?F�6CL]G9�^e>d+��:��/��@����@dU(
Vt1� �����'�	
K9R@�u���7����@����vMޣ�"P���M��������C��j�mG��|��B��'��H����k*|�Ї��y�s���Xы��kCz�7�!�t���=�[��	 ��h�m��S��R<VP��:�S�˭AB��k�$�(��W^˭��gU��_��#��U��QK��vU���z��q�v�N<�'T}_�m�(;K@�(=턠\�|}�:��2��~(Y1]l���^w�D ��]��fc�����+[��A}ϻ\�)zc�_燹d~i�×��Q�T��������\�ط�˪�Q.h��u��/��ʭxhrc� �J@B���i�054�BsT��᲍������*�̽(g������My���g ����Cc`��Q=�fe���(����z���O�i�ߩ���?l��_h�@f睪�������;����)�=��*[����}���`��}�{��~��b9�Mv"�zŪ&&�QR~B���$bB�j%zߙ.M���ѽ�[�e���a��ţ��l"���kh>�i`$�h�O��m�b��:d�]��{�Fe��A�f����.���q)��iz$	R�B�.�c�D1E�p��~E>&�{��b塂�p��&3����3�d��
�w/���iW�W��oQ�-�ʊ~���.(��u?[}ms�n���z ���F�M6=x�qh�I#���R�(0Q�K��cm��z;�͠���j�Ee��{�����n��ֈ�k�~5j�d�3����m�y?�6�o(@#!N�o�M��]^FJa,�O�  E^��p������~�S���s�,t#ltW��{�ч0�$���<���s���@~״ڇ3�4EV��j搲5:J��{�M����JF���>�[����ph #�AZ^0�zY�dP9?�{
Um{RT�IX �g#�D�%��U`��V��'m�n�_-П����.S�B��Z#�>U �'��a\+f��\�����r>�z1��K�������Ɍ>�жV��I����?�of,���*K1��y�J�&�ŕ˰�6ҥهD	㒗Q*8Q̨� p_,Uպ��#N1���l�(�힑���3����~�0d�F��X<�p:�,<��]+��N��We��Oӳ���Y\�/��E��)�\��XA6��JB��yc_��K������{�#&����L�or2R�So �Ȫ�	���ٙ�'���w�K��c",&Шh��3��L>�P���D��'\b�	�qӏ!�*y�a�w��a]�#�'=�~d_4Y|��z����  �l���}U�����p�HӜ�'c��?]N09�
���u}^ߋ�Ͼ��
\m�H�)�h�0OV��PH׻�4l���PO����؏g�ӆ��j�� +�'�du����:=��$��c��)ɯ�b6�lS�m{�Į��s�)���o��*؎Y�h:}CR�gL�W����4wQ�������@�h�NK��F�>Vti.�O3t}=����k.hv��L���^~|
�u�a��!<Y��y^N�G~��`�I�Q����|1aGb׶I�hNv��b� "	���Mrw4i�W�ie8w�ro��^Fߥ�>idl��,vŏӷ��^m��):B����v��2Ԉ2S�����d�'
�9z�G��>|`u���T)y�{��� �h����Z�y�BV�5�  {#�g� ������sc�f
(�󆀄�Ȳ�;L�=���=SS��u�Q���]�jnfQ	��a*oge����ㅱ�|�`�6��=$�w�ڻF���?\�I�$����Û�2���z���W��
�K��z�ﴸ�g6����YґS�H�+7�a�+�2n���7�E��f�c��I^l��6o!a���@��!\��� ���A�h������?��As]����y�^XIv,��BnlQ�4��y�6��\��J��˭��(�P
�UQ!:-��!�
��~	���@��帋���x@��l"sk����Y�ζ4 �:9��Ϛ���c�A�j('�qk�<+no�TP�p��$�'K��@��+)Z1�	
3��62�����[�!����oH�FG�u2�Z�GέЅ3����f�
�p�k�K���m�����i;Ք��KSfdJw�v��x���F��^F)(�eƧ��8�4���ms8�X��O�U������&��
�)ԍ�� 
W�W�{���-��"Tӓ�
1�9<h\�V��)�9�K��3������3��u���H-��G��r�C�t��K�[c�!���ܜƏ1��P��m��X�W�VW~�%(�C�l�d���	�9�����������LWZc��;����_��Z��;6���w\
�1?�d뙷( ��ߧ��V�6�d��]�J�-E��<	I�X���Z�u�8�Drִ�r��1�V�u��Z#��RJ��J�A�����HmH5q4��u�Ew.2@o���!#��Z;������Ie�Bw�X^X�!�Lj��`���@���\�/z�W�ك_��%����W)�rJ�-�w�����	R�J:��O�)��kpO�w"'_B�i�k*���l��t(h�-��kC�я����-�";W�b�pG�׈H�{~f�g�sA~�:Ih���G��pC��^D/��I���n�w�'��*W�B7�c���uJ���e�F��lz9l��cS"�M�Ȟ����]1�J��!`T����D�1�@{vG/��Ѐ� �s;i� ;<�6�^�����Uye��N��aUx)��S~f*%��k�8��V�Z~�+��Gk��XD��5u� �3�[��-t�T�\x!l�=�>� �MQ��?X�>����$/%�<���*�ބo��;��e~G<:z�r!������X�:�ǪN���%�����J�?�8��cH��{��aC�/�p�_z�� �X�8@����I~�g(Y�{�=>�f�}Cӫ�!��Y�?�d�%.&��E@e�}�Q����"P���R{#Q�ӎՆ����>ÆV��L1ȴ��L۹�}�L���b:�@[L��{�*�O�:HW H#�xj��ZY��<l{.�;���0ߕT��ޚ:�K}m��s�?RZOт��:ɇ�Q|߈M�5���@�G�o[��ڿ{��i\K��F��ZO��Ci]�/�![b��+�Yك���v���Y���)m��V�-WӱeS]o��n��}�.t�
���\a!|�*,z�ILn���Vf�[�AI� �{��������3F;�6���G�&�*j����7(l��%u�L$�b6��,IC��&D���b4qe_�7r��(z�7���ԂU �=�9�.̗��!�zn��p�3�K��40("��[n��+Ր�VE�?Y��奄�8ȧ�w����Y>>uS���ۡ®#;$����GK�m�4��x���5J���7I[�����a���qRj���� q���%�� ���] U$���Fi���o7��*�5�n\��)Npm��#��ݖ�7��1[�B��?��Byʆ��j*��x<�{���M:9��n�E�<'#f�G�q6Z��3Ƒ4��~z셀I��O��q���-�F��i�~�64�̥���e��2N.���Ů�!l�@��q�']�&�����6:s�����9��UgL�؟�s�T����d�ɂX^�sQG`4�#���2'u{�:���Fg�ͥ`ﶂ��Ũv�md��چ�i <Yc�����$�o>d6�>��ZɿX^�3EK��q�R+�&"�L��#�G��m�fL.]�B/�~�픩�\�x5v�*���򰫯!�>��U�$J1X�c,hb�ug��5n�I��zF��M�P�ٞ_Vg
�65�8cXx×��YO^n����`�2NK���z�ee��W��r,���=\���Aڥ^� �uC��(�^����CR�'���\N��U��d���=٠��$�oм��@�P��<e��w���.iDC��s�O$��HOVS�>F���U�t�-��*��aw$��`�/�<V����(�N��xB������eI�	Q���}L�@X��=�E�`���JK?�N���Sݓ�"�ڜcX�X���e~?�.��)^!Vm�����=����x�]?ܨ,�r`�_v�Ln�o�5%�Oo��z�=	���}���А�g�[S�ۈ�H#���{�y��]�W��s�eu�����v$����.ൄ��S9˴`���<�H8D�� ��*b��}n�>�lQ���w
�Օ���!��&�ÿG� �a�}��~l���XPt��M�����c��=��)�u �U��e�0�CΙ�8`��R|8G ?�{Ly0�i����FG�6��t~O���`�t� �BOL��f
�|g_�ri�Ŗ��+��������CA�S�J���O��h����M��(�d����>�Ɋ��"�M�j7��E�*`d�W	4���UȱU�G��o���<��Q���q�"?*JB/^e�F���4�p���X��,i�p���?�9Ņ����G�@)���^S�?58�m�4)��l]5�}����䠔��j��\Z�+}�Q}wN�<[��~�/��$�Ӛ}9�U��0�?^�
�B����j���yq|�����������ݯ��3{��H�G��{�/��pa {c�i��w-��D�6X��[�o�����@%.l 6���S�7Cm�KJ���5Ǌ��cr�k����Lz���↺G�����g؂���T���g��[�RE��S�/LO�-=ϔ/I�@���>T2��Ţ�/�V�����Y(�z�����tr?zo)z�%P�
$���w}�~O���aC!C42f���F���`%�&�з�X�5m��r>3��p��"�>*|/m���
����eϢ2�*��'�`����)V�,+�f
^9E�}^˸���@���7��KeM�4�*�t3)�0b�Yq�,B'��mE��20�0�R;X��~�I��{;��*>��O\a�83WB�H� 8�eDx�����.@>�`k̩j�Ɇ���U���a'A��q���$��VWv�y��|I��nz>��o��@�	��m���s	����2�n4A��.F����?\��0,�ܦ��*|�,��x�	v}� �=��޾��a/�����/���}��ddF�Z>����C�,@j�,z&G��`U�(��-����{c	tV͈�eSg����G-��V�?V`H����fG��߆���h�%�0p?3���*�ŗݱ?;�r�xω���c�R��4���7%�k��#/UC�r��K-�h<�;��3R]ƓM��yUyhX����H(��VbO?��3�S߫el.�X��-��3����,�Nw}�[�%P�^`Ez���
��ǭ�=" �*e�����Z$�P��u|ި�^-�"VOi�M��PB܃�LLJ�� �$�i�[m���3���i. !�LA���5�0-3q���c��j�JT�(ȼ��0��]D��T}����u��C��c��l��4A�+U�y4)�#��JoN��ɸb�36����;����7Je*5w�Ϭ"D9�m��R���2�������
�R�)u:vN��V��<-곢��b��(���6��K��$�O?�smP�V�Ɣ�Wb~(s�/s�T�:R�t�f�/5���ʕg��g�uh.�������8q�T��o��C�Ԁ�e�u]k�r����c�1��ӑ�~D�#o w)�\���c'�v��3����^�v�v�"N��|r�9JO��� (��{��hS�:c D�ç�u�%#Q/,.ֱ�� ������
q���fd���3��=�����x�DؐzO�>&���a����J��o�H��]d�d����R+e���z2���x�k���<�%�9��h.����yc*To�X�bhm���饆�N*���0��}��:
"�=��t����Ғؤ�mQb�هIY��jL9Kp������;�8ߊ�˶�ϵ�k�K���]�9Wt&�m�P�C1�[$�5�P�$�l��Y���8;�{�_�	�xq����(�*�����^}_����ZlZarDJ�ߖ�ñ;�=��K�$����Z����lV\�S���o�@0d��Q��%�,�έK��4y`��yN����-Gx��z���"�+���Ȣ\���G'P�e<�8����]h�=�-��)+�� 4���j�>{#��Ώ�š�ڸ�~(���u�~�������X��ۀ��"*VbxL#��7���?9HOLe(�#�����z+U��T����}���Ȉ����J;�y��7t��~����ñ�G嘔IWy���{?(껻b�E.�� �'�:-�I�Jy>I�������9Y�W�
��X�v��Ճ�0�(���Φ
�yE�c�/G>F�⛪|$�I�B�L�wf4��O��^��.3_m\ښI��^�&:Q��N����;"?">;b���f��91�<XGm�v���F����7�Kűܘ�FJ�zj-[�51��Н�z���%��ϯv�k�$g6�>�q����R�n@(/�\�#���҇��W;b�e"��ov�=�r셧�C����h�Ć\x�i��$�����+�R�c���Q�~�0~�<k➐3������G�:O�����	�8��H0O�.?!���'�������d��2� np�F����8S��;�R�^즻1������O������ړ�H���I��2��"�jLVoz�;�)*���z�7�=:\ea6�㣆}�9�λR4r ��RʃI(&dkP�bƬ�V��^��񊰚��fH�����؋���G��J�F��C~R����Z5�ׅ�5��{�\WE���5�?o-�^���W��g)t�Qi̮��P:N���������bu��I�x�A�C�#l~�VFqXO:QI[K�Ŏ<Ȣ���o �}"U*� =�C#u4>�#�=!����΂���:J:�-tDŜ�z���h�������:��	�R����lR�F<���2�at�_ �T�x���]oZ��Sá�;���\n {��u_�����//��{���H��n�}�d��X~����Ղ��Eъ!���n�=g�P$>+�Px�h	�
Χ�=����<�����_��E��Ξ���{ꪀ�_�Y�q
�w��x�[ymCvVn��Vz,pBӫ��Q���A+��Is�8c�����-`��tCE}B���85�B��fX�����b4"hnP�έU�R�'�;�[���)x?:�uT4�9��{��P��6on1�H���@���y!]�J4�~w�B��o�_*ష�̕�[�����dxK��XUwLp�g:B[Ht�VεzCEُ�MvXߏ�cn^'� %�Iy�1�v�A-CR��f#�V�䒞ۨ�juU��h(��6gF4����s��s�q�E@�-��d�����4;�?{9�G�^^�m�6�FKi��F�Mf�ߦ�5zd�듓����J�S F��
�@ϙrΚzn�m�H�p	�|�5%��uu�ddF��Q�	^]�O��s*{��z�L��Õ]�J�S�%����2-rd�Z~�Ħ˃a�r�q�����B�NZ�����K���ӧ����DPn?��,'��Ke�>�)Z^?ʫ�,�����y�u~"��[!�1�� �ˣ�v5>��O6��b
.��W!N�F%���Ҧ���GF��-�e�Z��B/�&��3f-�������(�F$�$��&��k}O�I`�}��7쩂�ڞ<TB�ʶd�.�I� ���{�w�S5�v\�2�8�ᙰ |8��3�92Se���=r8~��>lIA�$���Գcy<�)��x'��*�)�l���>�ż�r�����ô;����<�.w�h�f'��9�q��V����tnV�����
�T�%ko��h"#���]�*ު��Um�B�e����~N>a��F�w!�ȍ�}�����H�s(��p���)��W�x�b���^#ᦞݿ��mb��r�b��(Rmf��0��X��Y�z�!6=foQ����2���A?�U���b潅/du
��ZdYQ9��B��5��[��l:{��)2���P邭ѿ���<z`�:-��?���� ����:y�E�b���C^���{M�y8y\}I �$3�ѵ����t������ʝ���-�9�lWE��)�2z����S���	zS`e4-)/��p���Tæ�o�iT�M��>�Z�o"�>�>֫�y�+]��7�s��0Իq�Y~���P/�AYI��*>*���-���S�䵎ʙoa ���Üi�~Xp��}
-m@����b���Z�>�H��G4)��l�լ���ͧ�|f\��H�.�_q���N��|F� �'΂����(��_�)���!�)Ob�9?�F��A����&�g��J�Q+��"+��^�Sׂbd��:�f�g�����F���[�G�����D�Rx�>D�O�&K�W!�L`�Q�jϜ�%3`*��Xd^9N�<�-̳(J�^Y��H1 x�UJ�
��`��.`F!�.[���K��<�ړ������JE�Tɫ�lѩ�0�3t4�ߘ��ZY���y:z��G���s�芷�
���GN���a��<��p��)�[k�X�0�Ę]S���bCD�4N7�c���i�A=Z��$�aj��}q�W��C�� ���\iE��^Lmy6���.�gM�����)��>b^O�˅� �ԛ�tH|X��~j��s���F|�8�����,+�r��P�5j���BaZ�N{Z]����mY\u��)A@�'�(�]�A��ԶFZ��f=���4&�h֭,둚�0�t�"_���������L�	xr߫�s~���F�#��B����V�'1�JJ�N
u�E�ۿ�`��;V�ena'��Ӄ�n���ܜ�j�3����C��)�m�i�HUhr���XY�(�+�f!�y3�j����e.Z_�D'_�Ԑ�p�Y����|�/�g��{	�+
rXL/[I�3�Z��P`6�bUN���C;��۴��H�����z��
�!��,��Y_�`��_�N���&�v�b!�R��HŮr�P��vS��7b��嚸�#�jkݱ��ͥKa��<�J`�$�6ۖ��uه٠ދڷ1��[6��S[�/ �^c�EJ5ދ"��U�rv�~MNz�E�W��
���ދIQ�^T>	���qT$����v�n>/�z�!�N�����ƎA+ϼê������W���fO���4���[l��	5�4]���s������g�@}�`y{��w��VƯ�n&}�[���v��A�n����X%�A�f$��^�{^'�PT&����6��"`F�g]�������6hO��~of�/m��T��'��}���K!44��YL0���]�'%�K�o�Z�+ة85t��!B�]Y��`a��������N����$͚,L4;	*X=�+5p��B��ʌ���,�p�b�c"�Kqno߲҃��=��G�@���f~H��)$(ӧX|�؊Ŧ`��#?L܇���:�^�́��qǛ"� �(�1�� O�Dpht�3�n�0+����(�W^�&Y$�emY��t�r9��b�NԱ�z��Z��L���S��h�_�1|��E	��8�/�' ��\�$��t�Ab�����e�E,R_!�Y�H�_`F�� ���1�N�-qo	_�P���3���"��R�B���n`��:OV'�ri�%v�?�3�k�P��y��mAp�A�_n�T��ot|8r泤�C�b�δMl}Hq��m'�4��p�# Y�XsB��<��>~�a���?豍^:bk�����yb5T��K���^ͤ��AE�>y}��w�T{����
�T�?��v�����(�Gi����:�b�o�8�sZϗ�!�I��a~^Bm��=@�����0#w����.T�!��R����E�a�~��k)�ss���a�'�w&�n��:�zt�j]���MB��.u�,p��$�i2J�C+�'Z�d�a��~�MS4��V+v�h�cg�	���֖�`;��<%��T2���^ �o�CC?�����u3>��-�ЫyI�?���#|���(�*�J"LkK��2��X<_8\���Յ�g"b��)��w�_0 &|w�+@�?Ֆ� ���A��j��i�%� mA����:�^	Xehgۀӄ�;t�]�6���6�-��>�l�Ϻ���1hN��ݳ k��#�u �!��R�����_(+�b��|%��}<�n�P��f��#8%�����])@���us���S�`�:��%ԍpf?4(L\�t�]t·���M��G�ؚ�T0�:S�N@'"��������YM&�fժ1��G�F���ڦ_R3����<%�X�M_�߹GT��ͶS�,Y�P
?��/)Ap0�W��~��r5�xq��e�	����K��U�`���>�g��0L�^~�	�&�@2�uz�<���Bn�G0��������W�S�|����PM�Ӟt�������j�>��l8ǔ�x����X�n	Oķ���'�������t;k�ן8�š%y(C��m�j��Q�<X���)��Q��!%�MM[f���dSu��鸦�o]ӗC��-� oV��Hŵ(���x�`� x[�U1Y�������h��T	P��Sl�y�+�(�|F��G)��J��GB�HpqDs����}��I�z;����}��r(��0���	�\N�B��~��8R���5�v�NC�8�йUiY�V��#�EJ���=0�9[�.�J��~��9\]�ſ<��:Q�N����I	�W�*+ �"��g�7!t��8���S�dHCJ�D!G�e
�+@	�ʶ�jÙ�-SZ|�s������m�[q	�n �p������k�O��-]���O�&P6q�g5�9��_�Rc!(�=E�T�z=�`�߁��z߸D�Ìv�<>Ω��S� rC�o�t�g]�:�I��򱶠��筴����{��N�4&
�fn(������7�q�H���f�e�T��M@��c���0[���#�S�񤯝��͋�`���⻽��OI�QY�.�0��2�����|�'$�M�\�Q|��O�+;11a���d�?��3���W/w�^V��23�������o���u�C1�ڽ-K�㇯#5Lʠh��*B�$�q��	TW�Z���M-Y�(�1�p���"�ߗ`��Ϊ݂�to�4}�.9��1G�$n�l	sO�n����a8���p��ZNG�\�cK9,�Y`�NٌSGT��T�Q!m29�\?�f����%�Pka��@����	+��k/J���or:�˥U���c�e��!�bѼU�dSAv��j�8�Y���U�>�_J?��N��Ov\�+"N4x >�������-��G`_��u�5A���Ǵ� ,լ�r�|e����� �-�ɟ[�N��j�E���y�!��xt���3��{���I���.�*X����\�:}��P�����[b�
�����$!���r�0Hr_�1@cg\�\�1�x��@k�29����+|h5���wV�y��9

�^i����q�J��4��@���rGw�_u�pA�D  -����9�a��X�ƾ��y#�2;IM���Y!�w�la�ݰ���5�1����o�x�i����ў��*,%cA/����[4��(�m�<,���w|܇���p�Mz��6�Z&=�'�箮~�lU��t{nUE7�2�Y�a�B�0@�I� pp>��ɡy�q���]���-���02-Ҩ���`�	x��P�2��l\�]��QG�;�8�u�+���M�:&z����/2hJtq�z�2��|��T���;�Xh(s0�$)�2s8w�;,g$əYT�[~���ք�E�N�#��]Z���d�5cM����U4����VFQX��]�Q�?rSc=�	^z��p�x�D�tAn���E�D}�I ���-���Rm��ξ~n�0�}\��,�h�0^�J�%I�u����^��2̈́&v�ͻ�Z�Z�lf�N+t��G��گ�lt�'��`�gH��qn?�<��a���@2��?R�l�U3;�wgZ{w����{g�b�^��]rt�O��H8$͢�|4�G�֧C��`��
�y煍̅`�$��ۋ��=�u�Y�E�Hq��.��n�2�/��B�`�>�Ք�'w��i�0�%��mY*7����Hv�t�¦9�6��p����X�	SMܞ�����q��b��p��E�nۍ#���>�<��0��.S¦/c2z��.Kh�.��a�1��t{��/%9])�w��o�>D2n�̖W��i���ʻ6��Am&����K����^��|���fp��M!�#/n�bU�l�H:K?V��s���h��)Re����i����5M/T[��VV��T`i�z�328.Q�i����Q!�L�V;�j��Z%�r���F�H��l����}<�L5O���4-][���_<����w'�ܭ#y%\��G�`z|%�Px�qQ*az ~��|��\expB��t�����Q���/]�xv�aÙ4�8�!t�y��Mz�s�|.J�b"M�w6Ĵ:[�j�{�
7_iW��G��*�%�RA�_��-�-�}Ֆ̇E�	�R�����b'l�J!E�}��]!�F�);�%��4^���&�x�zjH���ŉ��U��'g��Vܨ���Z@�L�W>rmd?� �(��6�� Z�(`��Uz.�d8�]�8�b^�(�x�����7TT)!#J���!De�'R�A��n�CXh��f���j7��b`�N�^�$�~����[qb���0�p;� �
����S� �Uy�IZ��R�]��޲�o�̅�JA��=-[������H�����<�)�z��0�&>�]�Q2���މ�7�����"�6f��D�����a�gNlsqW �CI�)����T(���haSSF|5lJ�fsսw�,W{ W��H=�&+�ո'`�}2}`G��5Z�����'�w��TE}����:�.ƞ�� })'2DB樯4=x����g&֗_-U��qH��_YE���Ǿ�+��IUQCBe��k����F�߷4��s���؇Lʜ	�)�Ij[����r�[��4n���l6>6��[c Q���'��~���Þ�	���:a�d��'FJ�<r�����G�0��?��K������'`XM���")�C2���IB�I� �lY�	*�����*]/3����V5�g�q� ���|�j�/���7*�/��ހ��lųM�{C&#�| ��FXZS���)�1<dp����d�
���m�m�8��p�x�8�O�����Fh=(��Iԝ��pϫI��pK����A��h�e왻Ƽ�j��({<�w+��ܐ����x~�7y�^jG��c�	�7�K�~�;P��;�w�N����n�M@G&�Ĵ�H�1�(R+�ڒrȘ�#�#M�N�K���S�.2}}�lP'~f#C��C���J�ev
�!�`і����O�3
L*e��L!�
Q�+��!��[@�V�����@�ˬ��WF�O�Z�
�	�l=�|�ƕt�lQ�f!�|�0"��gX ��~��L>3�e*W��C]��]:��F�d��x�o��O���Ju+D��j?��
cBԸ�]z�H暠�>�����(��}�~�s��˭�j�rC�\��c�i�]P{�F�$G��;�t���s �r����-�����{= T��j���u�$Q)A��p�a�� �2�=N���I���(��-T_��b���KA�0�����_g�"I�O���;ڹLCO��o��@����3�Y%��hh^3�c��#����=�}���{���7D�<?"
]��pX�1�~�	^� �d$��Z�?K��6�m�8J�B$��D��|��d��w����� 	JmB�HV�+��Q��AV��������S�Wg��|�/��V`,D��|
�<����F2��~���UYt^ğE�n%��N\gۻb���:a�=��R[|��{�T�~e��ɧHY�m jD��/��wL1�-B�ɨ��h�#��Ua�+7wp�㡮�%�m;�=�)�5�
1��T9ɟ��WJ���:�h���[��J���!�9R���u�������a�c�\]�r��u�`4��x���ʻ�d�����X�g�Pϖ$�(d��˸.���{߮�:eq�fF���ǵ��&y�:�8��Hs+.��ֶ��\��zhS�a��2��uZ�A�Ǽ�$��+A�>�l6��4ZZ1醜�y$���#�)��<X��V2k]9r,5m���?���ƨ+� ��M���U�y5�Y���#dޤ�})�G�\��.`�ˤ��}�a�~�J�cA��4Kx{��9��<�D�'��U)F"�tL�="<q��Pm���#����z@u�d���gKZ*~d����Z��
Ot���6Ê;[FѶ��e��Ԍ��3�6�Hq<����ls�~лe�q�G�UT��(�wR�C�b�5|Wp9��y�`��"��c �-�>U2;3 ���� ܎� ��ʴ?q{<�)���"򙙘�+h{!�W��on�H��TM_Y�tюc�WJ�n��¥������&~�4�`�3y���8g���x�n`Q�B�Sq/4%� V>H>Y����g���)��m��a>g�=�p�?<�Ox;p��s�fh�?G�TWO'��2�9{�'��ՠ�,m"�څ=�2LӪ��c w����Kp��c�>H��J��s؆�������L��GW���)��qQ�ΊP2� ٧-�FnZ��Ȭ_�*��il���B�N�큚�JO���*�gJ%�	̯%�<^u=���r�%8+Ap�
'>Evs�qW!b"2��J�BLk�d=w��֨�_�����{<t�ح�	?MZb	��絿m�OdFI����#ፆ�>_����j��&j��ȜN�堽�n����c�|�"�G��j�FI+�"�f�������Ї@�H���k�����w�.z=��'���B���,�>8X*���e�ӴD�??��<[ߐq�+�5�x��=5f�p����������י�6D�8�7�D�QmdE����%��G�T@�Oϰ/"�5�6�	�8~�9����s�,� a����x����nk�
�����
�	3���]��da�k0j�Q�����5U=2[Y����'ta
�r�����!m:���n�)��ג������ѯ5���
�K�S��T��׀�K�GA�7Z�ή������$x<ۆE��p����)�y^��lu����\|Q�!$��'E������-!A�J��t*ݩ8(șɆ���5��%���.����0��p�����m��Y�����7/���B���2I�[�ŏ���Ӿ���	8
���4s������Ɔ���8���I�p#V-h��sJ�7�����:I%ms�2���PS90�:�XL�1��Y�8X�S�I���*c�D���pV�H���R�����7�t���<K�"e� �֪�U?��f�f��s�k<,���ȧ2"d���������8�~�8ǧ���x�7e�Iqݏ�9����/���}WA*Ԯޓ%���+��|p[��p��l�]~��!P����	�@#/��g�#E̟P��WaV�t�5pEz�*e�ɢ�+��ҥ9^���rCG$.�i6]�U��ҋ��{�[ܝp@�|����-ӆ�σqM��(8
�u�����¹��sTb�)�(y<�/P喱(P��Z��me> �g�|�מ�u%5\��.�p��	��a�M��n} ��JSj��J����y� {wۧi� f*��ƒ��O_�	�=uGv*���\ؚ��� c�<&p�� X6Oɥ�Aֻ������s��w>���D۰��4O�z���p�"V��|�0���әN�n��vݩ���pǐ>��Ɠ
y �T��f��IV�Ԑ/�q夘�}��n ��.Kl��}J���㿵�$nu�o�쎰��<}@�h��($a�&n��!�s9�-^��v�B�6�?�Y��R�D
(	���n-_Қ�Dͨ�`���sXWZ��*��J��m�X.b��dr�^��O�zL6��.1I�.��.%������vW�BswZm}�<肃����	���~>e]�뵫��g��j�	7VK��Q��o��qJv�
u:�
���k�,��v�z*,,�egt���{5��8��y���+�x�I�
��: $#����.
y����Q�����Ho6�=q���"����ߌΟߛ�/��� .$:%Cl��+�hny����?%��̪�j�G#��?���+�TkCF- u`�z�®�P&��U��;�羵��C'�?/� ks5�&T��c4><3��U�1@wۍ�A�(�Ah���)KpF�|=Z5��%�zWpM-X��:ʭy�4豖�*�B�z����d�l}�;�v����i�P6)7�BP�n��)}#�]{��5�M�*���Y*���.c�.��ݝhO;�U��pDV4�l(�l �B���x��$bw�{*`����[ϻ���攬�'*G��Sd+���7��r�_�h=T�/�H��S������i�o��?��@�j� Sy]��<�A������v��\���w�ɞ'N�����/�/�A7��0}-	̑d�(��"�K>�/]U�_3�$�6-��O��"�L�pF�]��]@8�7~�,�Hj-��?����+���غ��>�61�	V@�J�TҠ=ޛy���
�?:��4Y��Py����� �t����,����ˀ�|Np�a� I��Wsmyt΍��aZ�/��!��} �6�c�l�*�A@�47�`E��[8]r\�z�2Z�C�/Zt3�����1P-���{n�3d��<nh'�"b�)<�yv5�3u���_���#�N4�`��/o�j=&
�x,�BeVEൌ�?�oe�n��4���w�gZPM+�4���	��2ᚽ|5fw��v^���������L$��4�����@�K�(�M����"&4���η�u�g�h~{���86��'�90�l�G�}֞2S( O9s�rWp���E��7�o)�(7|nO(g����ާ�����燳�������,zyp�Ťݤ�l�x8�k�v�_�ժǶ�=^j�R�yw����K/t�Q��,bڱ���J��G9ǆY��@�4ٟ���?p+v��jo�M ߇5�U�	H3ޢ����c����>���2�1!G��["J�v�W+��F��ɕ��8m��1�j ��g9��Ay��q�l7eh�Y:I�ɊL� V����VCA�{[[�]�e?�t����v-]����U������KB�By�ۂ�{�W��w�+�.S��q�9B�z�NǑ^�2l\�l'���#�A�i�]���wi��kp�b0r��4�Ϩs�mD�v�����:����6L�o2���K�D��Ņ�����83���l���J��X��"�H�?DY���f��o����a���t�F�l�|b�iąIuoI��5�*�{�F�7M��[�&3ch�T��������M�h߀:;������{�\bê�Pn$��6��L3��s�bu��J�(�pn#n;Z����5�O����"���[O:�[}��3�4����z� �$"�fD�xsyw��(Z�4�u�M($ݻy�㘒wSd�#��e��yA�"����ͧ��}>���Uw��U�Չ5A=���Y�ل��yJU�s�0"q���4��}�v��w���%)(�6/��r:6���Ԗ)leo��K���aA�Gv����TIh� ��ߜ������ς�\/,U3Z�Mb>�� �$�#�'����~�ez 2�nh�`�o����V��q�C��M4��=>Cg��Ԩ�C����~=ʩ�����]0$� �z�NHsO�����֭q�9��-����\K�����U�
UV7����- |��`)cK����qïߍ���W��3����1�h���
캆h�������o�"�m�����r�Jj"2<ky\:�"���f�eW �Q�s�N�]]a8qޖek�t��F0��r���IS��_�փ��!8s�ٵ%���;���L� ��ٚ3� ���_ɫڥ�[ԁ�J�T�;���K��)A���nR"�%�� �u�~��^Ї̤5���ǖf�H�<n-Zm��[N]D w�Sn-�L1S����|)+�pLc|p�POǰ:�w�=ķ�K�E�[o��fښ�B�Sٱ��w��=��I䊫ģX(g>� �`��ϫ�`��,G����Tn�̠���Z�)���䋀dL��Wj��}�0�
���U f	�z;�C�{�g(�{~ٝ��!*E� ��f�-*y(*(��2)r6�[�N�/Z�����eW�-|��{�M|��"�`&o	���'P�q�u�wV�y�~��t{��A�+e�B�eS��{��3�Ј����+�֪���D�̂!�y��kf��Q|��ԁ�\#q�K�	�^5�uhTv���>ўY_1)9��B$���c~��l2T�Q�/�GGԱ���+)�q��#{cgS�h������E��0n+�R�n��##�s]�J�r�!����9��`� �Qh,�Sf�ϓ	�I�s�E�����`�Sʿ��<D/��A� �JՄ�ף�#�3�3�>��6O+0��;�KAF�5����Ĕ��ag���,▓�:O��a2�ݡ�|�q�w���8��2�Y0��n���VK�lϿӭ�ݗ�Ã���̈�P��g��
q+�6��Kq~
<�����,����U�o��GXY�	K�;�f��� #�ϊ6?��j����}O��^v��x���f�IƳ�ߣ.Qf�T��:á�x/dU�����\1Y�ޚp���}e5So��]�NC��Nҫ���Eۣ�s�M�xB

%}3�֣���|�I������O��N��.�����͢��B�=��U�uɏ�Ft:���wr!x.�p'�ePM��Z���>��GF��'��_s�1��S�����Ԫ�lw���/�K_�o\p|�a�Y�5�~�D\G�+��K�?�,��\�[�r����~1[,���)>���)�I�Jl�%��lS��{(� ��=4�(���\y�L,��&w|6���+C���A7�G�[T���������'�{��CX��7 E���\��Ś�Lý����S|���:|�}l�+���|Q��h�}�i��P}sт�پ�)K�ѵxYv|�1��.�����hl�gÆI��A
N��8��t�N8�I���y�X`w�3"���1`|���Ϯ)Z����zi�P �Ȣ����9X���x��x�V;;, ��=z��4~���Ȱ�`�`(�A�zh�r�+�̙J���1a�K��n0��7�_��Q̾|��p_�+����36���=Et�"`������%���C{�v������Zu�}7�0D��#�^(�y�v<aI��1�%�LW��J
pKv��*��i����@�b�J �eQ��?�Ыm�*k%�����a�3Q�&�f�La^;�s�_i�[d����7n��S� *�ub�Ԝ*� ��]
���~3|ŉ\N$�5c�7�륱��x��#X�SpW?&(M 7'S,rc(�{����,��߯��4�'���#�yR4Q�)��BYtR�_:wzw���B��jm8%p.MuS�zT+s>O�򜋴2���W?�7�Qz�=���G��+���K�f��2'���2�VƏ�5�ˍ����ƍ�K�m�����*9��)[�s�N��c�/��Wj�\��S}�)���^ͬ�����d�l�8D8�J#ņ���Ѵ��$�,��A�:e�$�L����JN�I�z�7�U�ZظI��Gl ���/��@Z�;��	��BK�E�G5W�h�*������1ޤL�pG���HJ�F+�8��]�Z(c�4��L��xX�t�k�/Ac;$fi��񊶜i$A�MN�fȶU9Ig�g�ߧ'6�o޶�mάj�X�"�eޞF�n(��R�	���5).w�:�]��Iq[�񛲦�#~�m��SG]l��q��dc$�tѽj�r���h��O�����-�ه����$4+>��h�,��S��[�굻��t��w)X3�耸���\㺌s7��Oe�"�7WDǧ��K�xi����1eON>�.@�7����� ��-	�9As{���z�4�G�$ ꢟ��Gqe</�)s� "��o	���'>���!�/�M��4yh`��Tj����V�H%r�U�9�}|@S��J�P������r6���bD��_B�{m6}��������~w:�:��Y�W���P0�� �j+���h� c�S����_j����2s��n��Ir����k�מaV����[�$�g�,w���;�,���^��eU5���l�i��
	z��@���3!�9ؑAfѝ|�e���/:
ݢU���zkrY��|�� �Z}�|^ �	����9;3Ȗ:0�.�כys��D ^���/�u�˴�i�X�!	vŜ���϶l�� �j���yޚ���� k|T�@�0��o��6 �q��_!���y��G$�Y��ձ��m�ʰ�1�%����;NX3� �/a��s�$�-����'/���<��f�S=��|^�kJ-I0~}�8��̺ ��Ұ$*��^X���-�m.,�i��M�.we��
cAʌ*�Ú*Fڔ7U�0�/1R��}	�'���ZD���o-�AY;���$È�29r�p�t3�=L�zv��X�-BQ0����\�	��k�H�[�߸�TZhN\&\��G Svp�����NCB�E�ዚ��,:!߃:u�ԅ�3J�}U��xmd��E4�XMtI鶳강�� �M;�&a�u����ы��5�0 ��$��	���	�w�12
��^P���?��J�6G �V���<ƛG%��n{%9Pz�r֬S>�7�2I�!Y��M�;buK�0��#������%񂆖��H��4�r$F\0�1�{�z��Cw�X��~G4��<�ߺ����_H��f��YS�� �x�o���>q���̪�dSu��*����RXP�GZKBF�F���}� =K���v��t��k��y�W�1n�Oq@7��X�+��O#A��1��S?8�2���w�(�X�R.�M��������k2��1ڰƃ��A���\�k�.zG�u>"���/kn��g�{w���o� �J��5����y|XG���ך��Y�>���u<�[%�����q��h�lv�)��F��g�ձ� �Z�=7AΨ�QȹN�����fO�CG��t�A�,у�X����Nae���j�we��m�+ƭ���uO�ŧd|IO�I+|#�-.��^H��f��ѽ�㒯��� ���E�!l�ǅi�\)]٨z�d�Ȏ_��]��͟*X�zR[��ȳ�R
���Z�?]�Rk���]�g�lx`�p��E��;��9�<o���k ���m��L�C7���6���GI�&Z�^�;ݘ�U�|bJĄi���v�tbj*����Рo)�q�[w���$��4��z#������o���8�N����$7�� w��b��8w�b�Ο�M"��� N����������f���;��Qi��/a�@딦Sr��\�v~wd'DY��x�% Rf����C��b;�Y�S
���jq��to�.V]?�N����X�-�R������(m�5���d��}��?e�P�ټ��U`)��g� �+K+�αJ��2�I���f�w]]��2QF-dІJ0O[ I�y�g7DK�>X\�d��j�6Hj�0:��	��j��çC��k視�l��w��x����Wl_Rl���y���!yTn�gK��[��;�=�r_����+.�3�Y�q���W<3R�\!6+'S!�������B������]h�K�
�F(���C��渢�|C���UB>�N����Ǡ�1M�j���;'�Ǚ�t�+G����!g��M�q��(e��rL	�%E7CMh�<��/D��*�4�w�L���52����Gdґ%i��́Q�^D�{[���zOV<��H�S$*�t UvbU��=���Nv�?c�3�I��a$2��~#"Z�;��\�r�x>��2ƥ�T����|%H�cw�y�d�U/�ӈ6��g3��j�u��[�� F,X���uQ�Y���&�:m�:s�j�0�SlԹ�D���4�l�yRл�l)��k�v$�w�x1�ƿ۩ah�\k���bu\㾖Qh���=ZהɅpD�eF���EgZ���F���ڐ��b��BBy�wG�΁�}c�u�Җ՚4M;����yL?�ÙF �t���K�8�뺩2`g��A� 	կ�o{
�̣DB7yK$����s�sW�[Y���O� ����y�`+�[���_�O] eI)i�]i�Px����Pm�˥�����Uy��
�<%ݑ��9��6Ӱq��wIF$a�����ȝ��g����ga�^Fk��đT�~y���e/�����b�!�=kˬ���G���6���
ﮜ�v�A����E������{l7)(���2"��~x-)k�X��4��5\d�?N��ș�r�?2�T�˒\���H�!h$_��o>]c2ò��y��g/�)֫+�agq���G?64�U�r�;���|������ʉc�M��B~�?Pb!�	>�i���*(}�i���Rs��*κ����#b�_��#rl��i9���:��ӉJ	�,ؖ�������*�8��x��4c��f��H���9��ѩ��W�^:q0���x��ꇸ�[��>���>��D/�@��J/$^��h?��ȭ�L~:f|�u%W��i�����P7�k9̴G�9
P�M���B���z��f<_��TfﴃfW�u�45cBrb9��A`͑�L�4 �UD�_8�՗�}���١�}:y��?tKv��Q)݁�v�7;'��Ø�6p��u�_�U���_4i�U�Nȁ^ �r�1� �^R��u����Ix��Cc����˕�{�y���Tշ�f7�s��9=����^1�w��H����`TՓ|�8_Qlͭ�V#j�4�#�Eu�h��Iy��U��l�������7��¢Q�e)�ܽ<w)u��Վup�פ����r�?�_�X!���`�W����9Ys���æ�.�E+�3\���0N<1��HB�Ba�F�]�sx�7`c�yQK�
�����Vg�}�@���xȜd�#*Ԟ)X �+���7��hh�:B��"�"�eU1� ��3�bc<�k�	���ĬCO�J��*u�;2�Ձ�	N���B>���4��ELE��?,cO�0{5�yEeR�Bs/����?�ab?�x�LN,8s��-�0v�7���%��H��Vd�}�1�#SF�����Ƈާ��D��~T6�����Ü��2#�X�R��s�z�Tƭ����`�w�G�{l��}8�mY��IC��|���I�Lō��t{�6�R�~.�X��*4BZ$��A�r� �~�x���6�d+�9^iV�p0q�s?�a�W�rQ�yT�c�'F1"}12�Hj-����%.=,�rx�O��O#{�F��ሗm�2?I�r���M�B ��iM��+�MY��]�-�Ļ�j��m���"����kFBj=[tvڧح�u��K�:S�U� #⺴���6���Ū��S��l��:ڧ�l�̾�$n�p�9n�'�{|y^>��/�*�R>d���ӯkT�h16h���P:�!D�M��˜�_�E�yu4�\[h����W�>)�vʯVL�Y`߱�p�Xi
���q�Ff䫍Y���F�\d��`�%�압}�.����b�n��&j<G?��,�"J�(a�ț���7�%Y�Z.DL��
�+a��>*�m���;e+�Ub1Vғ[�db��ǱS�����o���LcK�Im��ff�Y��Q�	�3� J$,*���a>a�hR�afe���E���_9]��H�L�uF�\Ş���Ӌ	��e��g�p�
��r��ﯫ~RA��K��\-b��)�V���j�i���8�&�BgxR������[3٬G�󫗐{{�P���Z7��R�^¹������3x�Q�&dԮ=���K ����y;�=�ޕF�at�S�r[�BZ:Z&-��P���f?�ǐ���Rg�v��p�z� ����k	�P����4�̏%^ ���M��׃�����W��5>(o���c�SY@X��4�����׳�x�,j�`m{�*����ٟ��� FGAH�3�H��2E/��[��?���U%�sdQ��]��(�a#�c��S�
�sU\2B��_��^���'zB�����
��7`N�d ��էi���1�-b���6ij��q�����|�C����D���Er�q5/����n�L���}�T�fל�ڦu�K&����<4�I`̖�N&9��B�[�!-��-�꣹B���vf%�3�>P�*�.s��
�����gb�#4b�.3��ڦ���c4 6�����S�a��{�3�m�9�Td�Y=43���uAR�>tq�c����fΐskg��]�B����"�~QDCѢM;Y����o���H3�����'��8"ļ%?�X`�	~�p���A&�������h�)\��� [|a��)�z���	�~B�����ܢ�%_�B����n��Օ2�E&���a{D�m���.섪��8����D3]�a�R���>wΨ��I�)H8��N\��런�pȀ�`h�h��&T� �ЯO3�M�\�}+��Y'�1�h��C��g��6�����HJ�E�l����jK��3#=�����O��q�7��2���:ru
h8���x���gg�Rۍ�-��/�����,96,�c>�����X�%�-���=��N�FM�y�'�ݳ���puR�@\�U�k9i6�;�h7�Oy�q��e��+����]�7$~���R��ڵ�2U��lE��N�C��U*��U%{(�7���%��Y�1%�LO �~�j(����,�©�v�l736����b:EI�a���^����H_�*�E�TE�vq��s�¶�.��F�(��Y:��-t�{>d{ǲ�U���k@f�7�@+V�y"�W`�^�Jډ*��r�)tܮ,&�>����/qPV��e��|@z��$��
�K��cn�d��� lU�9"�j2�q62Q=O�8
g|��{�!=-�JqQg$`�6�j�u���8X�-Ͷ�2����͵�)�$p�I*�2d
�@�R^ʫ���G��|�.X!�1�/h:�cB���HOЇ�ڨ�߆����Z�g+$����w��Ke��eY�:7F�f��Wo�v2�:,n�L��#P�9�%�x;�9�JwS)�Y�sg�0�%l9��@�=�G� .)�M�GJ���s*<|Oet��0Y�*'�^�6�Nj�C��܂t�iJ+�A��ɶ��@��ѧ,����ԻH�G�=�"�e��|��G����dJ���A�U������e�����F���d#5p�-^\5rďdӭF1x֮�$o������V�C�;�IG�BY��i��࣑28���sY���?�3����Lp܊o�X��U���R�D5:��U18izZ�=�_�������r����(#N�J"Aю���c�Z�ޕ�z��+�{�'L�=��-�p�@`��|&:���ڻڸ�{Yy͒�,�'�~rjk���so�ha1��Ok�4��?"����m��X�l�N%�PW�г3����Oe�5�8�+wx�Ɨ7�`�#<ވRi<�vu6�?��~��fXH��������n�\c�G�w��f�8�
�U*�A����=C���O��h�%���-:��A�h;0��<&�iǂ��W�M���u��OuLW�X�҅�FD�ruﶒ.�S}`�
�o9c��m�['(��j̷'�+[�G�L �w!q�4����ؗ��,���ٙ���J���d�� ��I�������ͪT1��� �&�x<R��(���7 Y��K��w7�6�����{Q�=B�>d�g����W7Ζ��j�X��+�j��d�{��ق_��,\G+:��4=����6 ?�%�]Aq�m-n��1����QbL^���TMz�.���o�V�:�z a{&I��G�ڡ^@aHO��#̅@9������ʸr�Ux�~��e䃒�2:FU3�W��aF����WX�/Cݜ��0�<��9|���O_c�kI���7ǣ�:�nS�W,�� ���&SB�`���y�g	��V���j��J�/Z�D �"򏬉6D:Sqź2�H�4,�tD0,�a�q{i8 ���u��0"%F�,tL�V�@� ��P�m�6�=~���Ȥ��q���
i��f._���F��ޙ��P��"hA`ٺ�`c�fD�]��T�>�o;���$	a�<���!��6���I���?Tb�
���;�!���� ��_��
��FT��;E&#�fڌ�*�H�4n�ߕS;�0��pr�V:s!\^�.�0gfо�u�����m��H��D�d��� 0�Ju�Y��������'CG��b��D5��ʪ�A�X \˯����5��/�Wu�0�7N��c{�)��O���^	���G�B�29�
��w<"��1���������[��I#�5������Hn�@��� � ƱԎ���/��8+ܾ���0�)��l�)�������(nl�́�(cT ��j'S�.$�bI�ˋ�%�2���!��NیVn�{ѥ���y'|�����{���=
�>���?���l�����ڵ����� ��S�ã�}���l��{s��\T�E�g�g�M��fG�$RW�I=xxʂ��.�L�VrY���!��o>~n+�������/b���_˸ʡè�C ���`=���z��kO/mJ���Q��3V��wG�y�r N�I��aɚ�+-0��9��%	8aM*�_#�W��ҋe�C�'5�lȝ_UIOe�f��q�'�D�x��Eqa�� 
���7x��f޻�G��VJ����i t�G�w2��;!����O�è"�t�\�>����>({o.eIhJ�[�R�����0d��� EqZ�E����g�E�~�2d��b�5���ʀ�V������uo�}U�^\��P��Yq,{&�o�p�Z�PP$�Л'�M�}a�
a:E��e �\�۱�L������oc$V��Y����C؋1�TU��B�ی��4����b��t5�u����ց(�����[��}�t����+��J���;��֣d>s���:&�����ӓp�/l��ֹ�J�9g �yBq��������)؝��5�%Ƣk|�i /8�B#������d��ݴ��T�z�P��#GHi,S��9�B���P�=0؆�h�e�0�!�޴�w�.���+9_��L�g�+��p��M+� �m������h����y@;�r%^d��Y��<��%%��O���DE��R��G���Qr�:k9�n�9�|�%)���<`��`?ڬa�|y|i7BSf�u����q��KGy2�-zd��|�+2]cѶ>&�`Z��zp�גb�.��d�
�*�	�{�5Ј(f�F�a�r�9z<�5~+Z����.�|��W�%HzD�(O�/r�
sϠ�w��e�S[ ɗ�حB��zU-<G�TͿ&�����Y~�v��Fy>�!�ٽs��@�0d�K|D���󵞧�*�J�5��3����&C��4&������G,4����[���t�TE�@m)�է/Sg��p�^\��sv����D
P�c(@ax+rG�̥a�"����i�\� ����r���U�3�S���K�:�1���G�u_���9�uG�:�U%&eh�%h��f��E�S�04�D����td��.JL�DW�c:�q9�e�n���3��dVLW]��<��4�7��p f zvo���S�ƪL�{�t���2���[�Q���B@L�hC9¼��jwVj�-�p�Ŕ� p��ꃉ�������.�[�sC�PԪ�������i��.�v��@Hy�L�\-����J������������ϫ&�x��J�?t�����t�c�#m[�?���9$}��gq��d�P�l��:����MM[�vR�B�Q�m�nM���l|m�S�TS�5ު2����#��0���,Ð�!�*b�Џ�V�@�@	E��X�V���_�H����<�`%�[�g����9�z����W�_;?����<�b�Li���^DAmz=S���0��^Q�7�8
��'~�Z�����VZ �'N����x!��Ч��mA8Xu�Є�D]
s����I��e)%)f�k0���}���~�����CZa�x��e�]��ң�.-�k	��'q9@�'X�m6��ӒϡЅ�:��ڛ�ݜ��5]�����K)]�[�&�d%�m��o�pzb�l�|�k�����?�ų�Q,�(ѯ��f���W5�ay�OR�s���=������b�[�bf���WGD���hL<�Ј��n��b�8k>ɉ	y�����H�j����sI�jZ��пZ�tXL�~��2�uD���Z��L�!��{E��3-g��V[tk���I��AC#]��1�dUG8����g��}��Óf�"�B�&�N/�VGK�d���x�R�1L`�R#Q��1ˍ�%��E��[5$`QQ�_���R����7 u5��w���ܰf��s E�Ԏ��/�xK�Ɨ�I���E>���o/��)A'�*�I��<����S�⢭WS��Q{j���4�yb�����H�?�#��?���$����ⵘ���ㆊ8��M[0+p��p�l�hr��(��y�rd���;Cx�,�,���kW���﹧�6��Q΢�����C~�k�G4�Fd� ��{��s�G�f
S�|��pe��4��[�ҽ�Hw3m�sq�`�J�Iʐ
�.�g&ˁ(�>`��W�B�}P(����{��k1�}�C���x䰋���#�G��ݜ��L�^�xV�ZX�gEl���(�����~&!��/�~ f����3&�םf��5�/D,�@8P]��Fƥ��}���J^=��F�P���)���?��Rp��s��Tu���0iYL +��//�f���@X��]:�l�3�X��^��$�Ϋ<���=;�����{T7�좒y������,A�"�78�h%��6��j7���/��Bp��C#UV.�C���NH��5_�����DR�j�&���a�����A�Մ�`������z�2OG�@���❏&�2��,BԱ��JԐY�	NR4��y�P�Ʒ��)�s�jt��[���xI��pMkG`q���,���H>,W|�~��Y4���A�T?H`��M�o͇MP<�N����x['����wyR�#Ip9!Hɭi��mȑX�M�J��ԥ��Zu�*}�y*'��=��>�0F���p��.�� �t��L|����ר̶�I�K��������CJu���[w<$�[Y�8��?�k�d٠�*���q��J@��s�1k���ʝ}�����n�?��+�'�6Z������h�Ȑ�껪G�1���A�,5;~˕��hH�q��&����7��Y_����������9��{vi��Q5���Ӽ��3��6�l�T���J��1ґ��ũέ!���L ����+����o\w$A�7I 2F`������c��Z|w��1�*��D'��&��k��#�,���������}S�����=�H�b�LD�"¤�PU����:0m�S�d�w��L?�͝�=H12���]�[��a-�ǚ|7�*�,�������_��)K��5}���3��v����Uy	��S������D`u�a�*�SE��S��Dr8x%u���S��N�ka���� b��K�mZ2�UZf�]��9B��U��Y��Uδ��q�@8��c��ࠠ�[�Q��)�\K����������o�$�u�8��'��P�y�P"�16c,�u�����!�g�X��⭪)�HDr�Y�"7��N���'�eW�R�2j�x�~k�ё�)�T~A���Ƀ����	s�Y�s�[� ��CNiYd��y,�i�]o�h1�1~��d�A��Ă��ݕ�T����$ �`HS��!��q��]�\x\T��t F�le��5�>��]��D��e-�u��szq��&*v�l�m���@�Q�O��&�Y��ƻ�M� �Dȡ7xx���������9$~�}�pg魏�p�],�&n�/�O*=ne�2C՗i��c����|Q9Ͱ�^W!������T.e��t�כթ��VM������)U��.{��H�4q��r���8ci�������pt���ӪF.�^������(��D�쐜�Z�ܡ\���v����%A��[��Q�\mt��fg`��]���9�{�}��I3�eb�*y\���
;QS݅u�Ŧ�Ҵ���0n_�X�3b���5&K��K�|IU8,�����R�L�*����-�S���ȑ��R��(.F�A֢6��q�O���#J���lf[�2:�Z��&6�d��_Āͣ����G���*,��<.��.%�c���kx��Ύ!.�v��.���,����g�|� ݉C/	�87��t�Vf�"��Mϝ3o�D
I�%ƻ�tKl�@�a��yl�phv��#Ei`B�u(���`�Cb6���ԯ�`��������mDaSZ�"�����k�j�|�9�⯢���� �;{�i h�+���82(˦�X��(B���*����߳-�%g+!ǁy%�*���P]�����,�Œ"�[��4�o�$1���~@��z8]8�ݿ?���IК�T�?/˞?�!�b���v����H���&�>L�|�h�G��[	�KG��X�t�tX�h([Ǚ��G{-UH�!M�>�b�q��OgV+��s��F�E^�5�@kB��}�*�&�X�NqK}S�!D�L�R[������7�������į{8V����</@����Id��mz\�{Co��l�R��� �&�*ط��q�b�����y���t�
��΁K+������F�o�23�>�[+��3���� ��%m9�f�Ns�!b�MD��޾��.�.�+�r�dd��M�g��\���i���1���4�EL��U���& �M�CoϦ��S2&0�w57�~���X<�O���M�H�J�펷`A�8����y	��q`*A��+�i����o���O?x}��.�\�/�7Β�uF�<9�6��i�4PQ2�SBUc�(��{_5m�F��q�F�I=�?��%�)^(�;�,6�7�Յ�S%�@�H�r���ZκC��l@���2�s�U	�ܒ? �� N�밦�١��-_��__#1z{PǬ���SI��^���<+���[��q���o2UW9/r`�Pb�_h��1�q�ѹ��q��ɕ3��I@ר��}�PS+vF����\�3P�7�m�W[�&��b���%�$r}+/\�삜�{��2b�/��6m�vIn�.�#�����D�Z-�lV����}�`�g���FeN<-�_0b�v����U5�B�$-g�ṷ��}Ӱ�Z��P{ڈ����0:8q6��"I}���C�`�F}韃�N2�u��FX�\��+�%������w�>��.��q9�^]o.4��J|ji,�g�)�Է�O|��ho�zP߸G�b�.UW�<2p7<�s3j�_��Z��R�S��q_�wv��{���5Lo��{IZ�w.��
���9�BE���G��	�ˢ����g�n9u"(J�S�&�����a?9�j�OwZ���YO.� ��=|X�Y���S�E��(y��� �o�ƍ&�k_fZ̃թ�"�����3@
4j�*�^��a�Zd�1��/��n6��c%`�^JJ�l���c���x)�@��"s:�ֿ����ߩ�I,1���S�����|����eC
F�l��VJ��cy���zC�4+O6�ቺ��j�sR��#��B��.(-�c��~�ﰗc��O�j�*X	�ɥ&�(>�im>:�i�>�����f ����t��kLW����n
C]i����{�)��&�pB�H�ˑw��<v��JB��<�[�5�9qk<�_�����
"c9w�'!q�tW�ɽ:�Tu�5��\;����ɞ�~���KC��Q�����rW^V��'����-���D��=� pG�ʾ��Zn R�]�^A@�hP3A������󯉳s���Ax3(���.oa����l���S��4t�����paPz�D��Ґ�
���U�%�q�l$����	�H����^l(�� ��O��Vִ��aN���\��p�\����:�߫��Z6� ��>��N_`S|s$�����Pā2��ȟ	?�	���h����*�{�'X�M�$k��Lk��S�%u]�$�`��J�X, e1Q"��桊�O��Ly�^B4pA>��,Mg�#p�2V�4^L5Ǹ䡒 �]$�-�h�Le�uWʽ��Dh\m��N��U$�3��L���!<Cn)�y��S ����˔;� �Z�T���k���"��3�+Δбu��:��L��,�����&Q�!J�e��5,����pm}�1�����) �߽jV�m����x#GxӼ�?F���	�B��Wq�߆Զ�l0��AL�=�0̺I+F?���Aui_��ڪ���[T	��d{e�]�e�l4H��&�̣�
��X��O!�^������+#%)��C`����RTH�W��kdV1ٽTψN9�&U
�W^��"q�`JG�Q�w�V)����]�&ͅ�92!'񟌕nV���R:�h�L��˂q�� ��)��r?���2Dt#"��nF�X*i�-�Y,8�
(��?�y�H�]i)E��X@���t�`�̸�TT�D�U�/gI�)/M�!�TCe_a�F��u��;i�)��,�E�_��ى�9%4�P��8nn� ��MJ�*y���HR돒R�@\}�G����M�AT�`���MF�f�Dc��]N�	��Ew��^c�d2���09 �O�� |Њ���a���ދ�:}Z���L:}@�����9K�����F�.}5Tw ��NY���c��K%J��ϿM8H�DIz�����0a�ݹ����v���r�Q}�n\+7�j��Sɲm��by�lw���{�s�hZR:b���u*�2q�����-����}g'�[�nZ	������V���C��b@nx�$�w���,���'�uc���')��V���ʠg9��Q�d�5�����
e��=���W!Eڙ�v�>����ΆZz��ґ2�9�����w�.^��e� պq}�s��ب*��Š��7?���ġ�*��������֫�L�<Ƙ�Ǖ�Q��Fǭɂ_#`Ͽ֩f��O��<ç�8��51�QE]<^�NBפ8���K�BP�	��@����*��ig��`� �R��s�3�-���ޞ�%��9H	���He��V�|�G*�r�<�g7�������B���v�cn	��B ��"Z�'.h-�� ��;�tIu5�py��p��{��!R�q�9�)��tH-��S�RR&��+�(�px���񉀙$�U�>��$Ըɶ��^\��<t�V�H���@���1����5��y�3�k����z�Bg�H�	#��T����Gڳ���WZ�V�p ���=r���7ݹJA��A�;_K�h�y��!,��;W7��d�� S������@����f��UG1��ᆴ�v>ӷ��F-������M�԰k$H��+���0�n��:��	%Ǎ!�c���9yTjȫE�(�Un�H	��@b��5����G�c[X�u#����[Gt�>�����\tе.�5������zz����%����7���v�!8Ԛq@�k�M���4�6[��}h�b+ri�I�����4�g��a��/}�����U�B�4�:v�'�rlf��k�=���|�TX�Ò�!K�\9/y&B;���,��K�9W{��Z����f"����Y���I&�h�eu��_�:���ңZ�
%����wN�)����>��urCvX�����2��{`��E=:���#�B���Ug�AM�K�s>[˪��|"?>�<��ظY�v�th��	շ$��Z ��A���x��B�뱁ꯪ��B�����'�}<�]�pH�u����~Ɵ6�>9��u5p�fY˸!O�8���f�'�i��)^,�-���KR�V�WЭV�5�CG�;��S�8�C>��(�W�%f˙�b�>�N�3�X1�ݧ�-+�$�p3x5\*���F�l��w���jH �N�4�Q}�a�g����t��n㕏��M}�#Hh���::��'K�j�V*z��D�y�L-�>!Na(�^�>���:t�jQ���+�F۵
}���ҕ�	��3�F��C?���L�ۈai�fh���I2/��0[#F��}]r#��@*�Y�,��� ./a?�t`"Q��ߝ���ʌGxr�������{�37��	�(�����V��IY����B �8#F��}ʳm�&�}�;]x�gȁ��+�p�zɰ�\�]�p�C*.�ΎKS�c+�����L`���t^�I�{���g5���+����JG�@ʬ��;2U��^=�;Y"��>�om	w 4��`̙��4���ZG��=��!W|�~ᛞ�	3������{��T��$�d�.�l���(�i{��3寕�@׃�'X��: 4jIV�ǽ��uRV��+�i�t�' �f�<�l+��g�Fcq��,������p�	��ʜ��uE_�W�fAlIe���l�˵r�/q�"��C������|�6(Zd�dj�B��@{[���Eo&�D��I����hvW���^��ԅ+o����o�3�<���*V�1�i�����c��Y�O�c%�?r��x������b��ݶ#�F����GM՗�e��Z][��k�o�����?+n�����wKR�@=���l#g����r��g]�,*Tx�a�ڊy`F�6�N��W�4�� �ñHĽӉ��NK㺩_�Z{��i�\��9��yQe���<AYY75L]����Zwu�t�؊x���{D��Q���_�\�B��B.��Ȑ��^�vϥ~Ԇ�+M���b�H��V{�I�N�L;��ߎpL��h�����֧I�"01)&U���}ڮ5���׮�F���حde��Ǔ��nv�����@��i3�]�Q�2s�2/Yqꨌ(ҩB�/��N�5��4mN�%/]�Rw���Jg�a�C�h�D1��G�߹���B�H�@ٳ�">ċ<�o�y=bJ�?+�h|�w������9��9�UmS�d��%��h׉�U�L�;~ܦq`?�ϫ�?۷{$!��� 積NE\���L"Y������c�p�����U�S�"Cۉ�\<U�'Q]�����۲�A���s��_mn��<�A�H/��b"��9�	�^��qG�2^o�m�Ix/C���31R:��x���)KaJ�g�4zu�(�*�82�7J(�'~H��خ��+������:쿚$d`������3�{t�݆�K���s����jƨ%��P_��pA�#k�҄��$Yyv���%�XY�<sǢ��'D�F�N��H�����>c/<���q\7�0��&�B�#t�wkc����X~�����r/�x��j�ҹ�G��G7ף3��~�+�4>��V1r�^t��ɦR �Ğ�EՐ��O?Q�ǀq�Ε�a�P�sB5�E-��-s��A�2�}��h��$���y�7���;�d���V��G���[�8�D��D,ՙ�P[�voXO��Q�WG��~�����7'{��)��X&њ>�~�����ܓ�= e���,áV"j��Vʌ���˘"��y����+S�b[c���e�Q	�M!�k����E��0"����+�\fLd��7���"���-!\�'���TU�07G��v��c�w<"�:mP|����Tv4M�����[����'�G��d���[j��u��s�
�&����{|z��;+~�R�/ζR;�1�+j���w�m��k�4�HSȄ������#�[�Ծ�����a�e6+W�0����!�;vqԾ9�|j�L<�Q��~Y9ED�%������z�S$\�fzY�6qQ�3����e��=4���Pb��PF���c='Y}聹��/D'G澜��f�)�Υ<T���;�<�M+c|����络���\��t�*��7�F��Lߗ�;5���J����EۥSF��ǘ��~*�?])��?���چh��x���Y;QG\����5'�=qA�P
ǚ1��,��ׂ��1,���2C%�}0�X#A��2�#Wxe�m"��ծCV��F���ۙ�*L��'4h��8��"k4�`�#7�de`�=U
�2 ٙ����4�p��co��:��}��h�e۟9��l�b�(�K70����k�b	ā��#�]�A�_����[ț '�wo�H�ֽ�mQ�����:�*��\G�X�ח��8 �����y�3��>S��Lt4��~gC���.�zi�V����d���7v�ϟ��?땭`�$H����B��Ď#��J]��Q��M��r�\�U<1�]ZV7WX�%`g�)�}��MN��򹅪7�*�`Q�ra߸��Ī���>9/��{$8�/���C�8HO�H�<�D}S��4���f����;�7%-D�=H�����CE�#
����RHq�NU�p������b(M�6W�?���u0\5Ɓ!c����/!�L��Ӻ2��d�,���_�4����](��+�;X�N�%+,)�e�)hS�.�i�BM���8ܘ��u��J�i`;!cwӡebRqc�v��$j��ڽ�_%<N�-�@�yn ݸiri�вW�X�n[Q*8S�����E�W'��'���@�\�T�t?�$[�h2	l���K ��*�q=G�nTQ�jx��D1�͸Y>��3�� �GV����zi[c��+�q��W�������|q?�楓�!It����̆Ωv-�<�
��Fy�U�CH��.�a%�viZR)o���9�+Px�LVф����@�7c�-d�[2'jf;���X�V8�.Q-<cc��R�h����������Gk�R�sĶ����h���R>>:7�W߃�5����$"�ţ\�ocxN�od Q$�w=�*+����Qs��d�_��{����ȥZ x���tWU�i�Ũ�hL�����)�U9(��#��!y�X#H$�E:uP�/����{�m��e���n�"����e#�9L���R��pf���,��F?�ۉ�c랮�:
��'�n�y���p/F-H�te�ۭx��8� �B���cgD^5�L�&OT����){�%[bp}<�5ق��I5�L��s�e�4G��!�q���l	�x�Aj�v���}+��Z�Ύ����g�@��FPF�xc��=w�J^(aյf�d�j����v��gQpۄ��k���a# ���'�{�h�j.7���n���</?�ٿ�$;<HE��1*����|�-�y��=�x���s��)3:~����&�<�/�`��^�b����m�mu��s%����^�0UF���b� �gz�$�^��1�����ْ�kD�h%�P��zl���ب�� ��\k���܀S]�Jp`):���.��G{KVv���ggg�ϥ��]��,������J������;F���ع�V���^�j�e�rBԡ�LsNI@����Ž� ���_��JP��{S�V,��
@ϩ�l�Z4�A7�s�;�sr@� L��ͯ;GS����\�nȚ�����>պ�����Z��wێ��G[U��^�j)1������g���%3��$	�r9�q�Ζ�7?O��^�4��@� �$ar�X���0��=��u^�wt���+�;&�άq����G��I�X�K��}�~�����W���'����a� �k��B�{Gxܕ�Ir8f),Ѽګf6��I����O7CT3j#`(Rz|*��V0�lʈ����s����:����Қ��D�7��Ȣj���u�f�ێ;l��2gj0D�=)KN��W�{VP�iu�H0ɀ����ߠg};�lʳM Y�:��:��a-�2��#�v��Th<�? Y��o�ۆ���)���qW��e�E*ӈ5��f=����ō�My�c�jٌ8K�0,�qIyce71&�*�d�N�����8�g���Ϯ�<��B�,��yo���!���:��Ku��yY�%�!F����@�L�H�l��Fd���t��:��`s%`���}�Z�Y�L��-�����/w?�V���s��B~^Ӗ���U�vt�N$J{ %�ʂش��\2�奊 �.U�=:%�����y�3%!c|ɊO�a~��.*������B�9�l{��{+餼,��R`��Mܝ��0K�T`o���%�ni�q�y�|Í�j��n��֘�p��8���L�!��G=�kҽ1�$��갟Wt��F�r��tR+�WZgTa��%+~�-ޟ+#}sr̜��sU��`dXw"Y�μP#��fѵ�[گ�ڒ]�@e�H�z��Q1��X�oi"� Գ�GX�Q�jn>���;\OǨ���xJ�5nt~����>,?{�fx*��X�5��U���B �0�h���\l=���=�Rv��2?_��w�B�G�ر͠���+_q�����9���$�Xi��hd�7��z/���H���J�G�4w��b%�i�BC�[0�,�M=�7�=؀5�����Vh5�D'��.��Y^W�Y������6B�F�H���I�|\���\�����'	����!VϞڣ���du��-J��&oԢ�z���e3����x�,���*?D��	b1�eǯ-�O��r��Ό�	��� wf�����?D��4YDl�F>�*V���+�d�mH�����D����ݼo]ef������$5�)%�C�5ރ!Y�ȯ� %!_9�G5�ąЍ�ǽ6�1��yV��`r�f�I�@n�ro��UH��>��&R�f���PЈ�ǘRA˾�ڌ�����]�
�C�<�s�z@Fʖ���9�T�#ު�����	�PK��ׁ�si�df��� 9��iH�	�{W5�M]��w*csaI2���.������">S�����>�!'��X]npi�o���]ܸ������M�d��^sJJ��3fX���lE�7�{+Kz�v��MB��&�7O}�i�A����C��ܩ�PI�Ϗ'c���f6u�[�)���1XF�ݱM<�IliB��b��6x�_���Pw^���[;/x� �7X�=�qp�8�K�Z�dl�ڏP�Dt���R��i�|���2��	�l��پ鲗��ԱSw��d��#��]\P<i~
1��D�U����-7�=�n��"S5�F ua
F~��l�K2�z��FR��C"�WܦC���&Ue}/a۹I6�-��˘^�Te��Q��I�M�W�������
�����9T-�FB/��@5��#����s���I�V�n�oSQ\��s�q���)��c�'����u���:T���Z�V�mm&���D��E�t=G��������sv��c���K�1s��j�RG#R�8�V������SP��]����KL��?7 G��kN*H�,}�G3�lU)7PǗ)դGȪU>��1��He��K�cKG���'��$��F�Oз�b�"s�y{�dM �=&I�#�tɼ��;0�`��޹���6�5�zi�:����9}�`�%q������ϑ1P�{7qh�u��CR�MG�j�9-\����8.��؈�ªGD�|̌DS؜�a�+]|P�!z�q,+p�/��<�T���U�l��xK7~�:��ͱ�`�M� {��~�~ѥG����8���x�?Њ��P�6��j�|��f������NN��RDsPx�{��h��y;�UȊM��'^�.7QC!�DD��8�1 ������!0!�xr�7L��]fG��p��B�J��<��P����x��݄�hGd�wx�m9�®p�Z����I����n%
��U��iWw�q��_qz47��\_yn�Ze]��y��R�ql�-�*D��%���Y�� 
�x���{%a�mn`!z�.��*��$`���9M����+z�ڲ�уÅ)+���j+��^��N57�,TA0.�������c[�zx�B�9@��P�?�w�V3�umC0U�W/H����RoF�-�g�\�4�ۯ8��TP�Q욙�p
v��6���^?L�A~B;����}�a �{8�
���J�,�_�!�	�	�d~�h�G,x\`"�*�H����b��0C嗃�4f	�ny��=y;���]��ȫg���N?
ױ�y"�t��Z^e>+=l@5���78����iC�Э��<�]ب�h����XH~*����I���r�dgSo��%w�o_J
  a�`�PU��U7�C�)P!@�#$)YP�3^�[E].�a���b������Tt��wu��sJ���DB3k�6�$���1 e"E�<J�����a>�����G)X�n�D��)\ҁ�'b|���Jݛ�w�~����E��c̢�7X��f��+� �W">J��C����u98ZA���F�0`#�f#x�7'��M�Ɯ`��1�������lt���lA�����N3�������iP�>0�u�v3��Ҫ���?'�9�U��z�7�����^��h2y�3�c�L9��H��zq�ㆷ�mK�1�y��6$�o��J���+-t6ئ�J�O��ݜ��9R�)4�����j>�{��x�SU�~�Kcx�;�F1�B
���P'����D	-�=<U$�y�	����#E��t����7|y�3���$��ކynR!�2�!�d�
,�J`�
�D���I)�fd;�	�w��9$0�KS��v�a	�^(@]�EA5?Y�+���T��6�2>~�3W�-܇.��N֞%����C>��"��ݸu����j.V�^�'��l�	�&�0�[� ̻b�O�9�:�����t##Jb.~�����1��Q !�%~�#�=勦H�m�cZD�ȅ�͝��\Q�Ĳ<؈9�/�<�=E��g�,<%�r=�2j+��-H��`���a>���~���&�v�'?��0A����˔+�m��C!l�3S�&�(��	!BC��<xnȱ`n�,��|I��*/��&��4z_$���
��v�:�[P��F�J�����y~�߭]Gg�R"5�y�YG�t�)$����4]#�sг��C�����ƙX��x��%*����Ąg��Q_9�8-����n���X>b�I��A�:/Ϟ�=xREct�[�x@e� ֆ-Kk"�X�����G9ȴ!�G��1iju�b�Ř�]��j�x�E�������H��OA��T���)��D6��n��3�݂��M��ǔDzS�3�)�G�D��2(Xj���\�>����E�Ǭ��=;���������p���ل��O�p /4PN�m���s爬��K����j�G�Lr�_��9{쏜=��0�]�8�������^^ڢ�O��hL��$���S��b3���D�Ub��V~��*8���^�-�_��풋i>�bѱ^I�S3�Qe�n���*�+�S�^nU�vVe�sc�Egbh�/C"V-=��Α�(wS�
��v�_����5��D�p��
u	@�F���z�6�q�#ZP幾����l��x���1��D��kv�G9�:|6RC���Cj��=������J�d��]E�K�a�x���{8�e�X����ka������>8�i��7����%PTa�/����B�t�����hx_�ڂ�)�;;��9�1���j�$�ӢU�w8�!��")!j?	cȤ�Qc0͛q�� �� @[�"�͗#5��!},�h��(�v�� �nIQf8(�Zs��'�t�Iֻ�4�C�}��3C�Bxhy}}lI&�}�r��`�8Ĩ�Z9]�olNR.��`Z)e���迣�M,Wt!�v�*C�mF`� <��\>�<��秾��_r><(��F�|���`!�$1ԍ�b�x⊂"���K��`�0�Q�Mߵ�J^w��c����I��u����Ł��
t�u����p��@�1��@ !J%�ES�K����4�Pĺ渞�;A�.�٪���	'�,NJzR܂h���ai5�!�ʑi�i�yU<�$�*���/Gq|�ء}�m�o�`�f��`�:�t6�6�H�%��A����z�灟���"���8S�� T_�P�� ��:@��W 6��{�u�����U�Q=� ����:_A0��0��5>?�~ӿ���;�$�eO���%� ��o�Q��10�����K��ZPiC�b����SM��`���W*�Z+��+�xE�av����o����v�u��@`�e��8[���vl���~��n+�$�3ٕ���I,�Tܣ D`f�U�@�m���i�{g8@�I�(��C��vj�b�1[E�����uc����%4�Њ�_Z���k}	�U��\urVχP�t���z�`3Y@��@%��eȊ�(Q�Rv��٬q��W���L�2k��Ăaee���%@�ڹD} j1c2<ծ�@���<D���@�+g�kl"E�Z&ЉƼ�;����m"����D����܄��Ϻ��>�/!�V9�2�I�7j�[����wg�νݯ7��M���JOy���9���/�Qs��|۳`���sb\u�ceٕDM&E�fڂ^d�~{�|d�U2�-����j�bz���0��� (n���Y|�����O�~z'������\l�]�Ai�] �pg��m���&���ܼ\"$�t,�g��q�s�ΛVB�����%8�B�B�~����^�%�z�#aw�i9V2���'H�����z~-T�#�S<�&��B1F�Z���d�ڊ?+_�@�''����E	�C}(�s���f�1�.��x0@�`}de~�����]��T7��c҆�_��y���2-M�q;��՘��g*�4�Kſ?��3�x��l5��Q\�P�@:?��S���I� ��p���ō7<s�w��IU7��#J�����|-��{�Ӹ%Iv��K�X�ö�J�2�x��3�W�GxBr���u���N��-�Q)W�muM����F��D��0�4̴c��W�/���O`����Q�ɯ���`���z��V�|����]y�Y��~��2��&�6~�	z������o���w��	��`��1�@�_+O���.a�7�4�n���^�����P<�K>v�ׂ���VC�
�����js�%Lkĕ�.YC���Q6���F{�AVg@n|Z��"=�օ �� f��t���PB(�ޅG<L��iI���&�5���DH_~���H� ��۵I��.��8������Ū=tz���uja�Յ^%�b��%t��ͪ_�PI�H�x@���콄G������˻6��v����L����
ZS��M��+����=O�pY��3�����g�u8�۩��H��{ ���aqK���7/�T�#p=����4�n`�c�&��0��ؔ&�tn����K��M����`��\zk�ɧ6ч�9�@XN���B�À0��Zl�Hй����� �T恸ni�V�v�ǹY��~�F�fkD=`���>�W��!�h\!�<a��aj�+ae����\j�l��+w=Ҩ]���P>�AΊh��:U0.�^�q�E��bz���0��� ��g��H��x�p��l��f�1+�����z�� ����mr���\x�:o	x��L��:��n��^+䧂70�kX���M�('��F��~㟕Xj��Z�)~eg&�
���#�C�.:5������k	�p%�b���}�<�P�y���)n@��G��������ȅn�e��gg�����2n��r�M�9��k}�V���֫��S�N�{]Ť�d⧭3%�rM����0w�SN+���1`կ�O���Z� �8[�`a�E_����M��px����Ǒr��$!�=1�@��ɜ�t�HFl�K��lE2���L��`�*uh8B$�s�Q�*.'��y��zs���'�U�_A��<�b�E��[�62�mֿ�v� ֋��l�ԭ��ZC؉/�&�ԚҫP=6]����~��y�z��4M��r��WB�6�G�bx��<v�7)�z>-�5�]B6۷pmFA���r�F�
&��`�)�4eÔeVBL>a�h�ߔ֑1��V�o̚��P����ߊ�-�<8�Hjf�H�����=ļ� ��l�?�r�C~�����%3���j�����	降q଺�Tr������zg�e3o���^o,uBj��0+ȏ���7L�U$��� �P�e|������b]��D	��:+���Vzi���u�7��	W��f��s�J��h�E��=>J�0@�AǍ7�W}W0�m�/�~�hO��$�'_�S+7���X�[x
7l���{�>OU�*�U9�N��?��1]8PUPȢs^SJ��.�7�R�����dl��t�?����4�q"3�I��۞�@ۨ��f�����.)���t�--/L~�k�G�M)qK�V�eR;7��;������LH�o]3ʼU�<��@�|�f]��1�K���Ӈ4M%���S�zI����ɷ�u(q��s�<fNz��t�4�%@�V,�M�f��h�)`(�`F9�QB�Y^�p����L�t�܍�
�{���$Yc��U��W4!�����6Q��ykǨј��Ϥ�����r&^B��q�f�����`=��������|�%�:Q�L���O��.&�����VR�9��6R����,/'�c�9�l��J�Fl�����ơ}v
樁џ"���`��B���Ji�B0���^��}=3`p�;㼛�Q-��H�X�o7�N�ҕ)e�?G| �����ag8C�G���&�R��7Z���wa]�y�z(�X��/�9��U�_]�>;�id+3�SI6��M�{�6�@3&���Z�}*��|�]ʘiaN�zũj��o�exd���$W4�X�7S��ܓ���(��b�we��8������8��[,����e Nü��Ԁ1�!Y�״����1����A|M@���ץ,�&_�f@�������ۖA�6� J���em������׶1�&�okPbj��
PJ~����n{f]g �g�Bz�;��}"Ț�ľE�gK��M�MA����)!�1S�L���I���0�C�)|�Z�}�n`Oo��d�k��%}'��;�cm�H}���\�ph`�d�Oa���o?��.QqU;��3E ��(M{a:�Ӧ�u��%���F�늩UK(?<֮C������`%\2��a�i='�1\�����w|��k�\��2(
}_��
�]�^T!e`��g�#��AI2��tJ0�i)�/e0
"����b�V~y_��]�6֠6[7�Y��
���D��0��ٚQ�<�}�Y,o#����s|�C��AÀm�2�Bl��g��v��T�"C��x���.F�
���
��y����ص�&N�a���;��!��t�8����6�O�a�?��M����ץK�@�
�5tO��ϢSHF-�喐��Kj��.�}��WŐ�\���0��9Ⱥ���$�eh��`z��6�!�:�w�G%�4�<A���33D��?8��+�����j�� �Q>[~�����vL����]��;k0���z
�K����H��}����6�z��������&o��it�6l��R�VU�;������g�n-0QPYIj"U6��J�&%%t�Y��� ���"f�]��_�e�ź�zEŃ�5�-�>����1&�H�C����}ƨ���6c&pI6c]�W���,�UR�N�c�Ɏ�W�`�2�������7<
Rk/�x`>y"K^�9稙e��P&�/'�������W��W[Q^���YU��~�U���׿�n�>A%x�p�kmF�=� 'W;�g�k����\`��F���i����i�Tژ~�#B���-i����\�\
��R���[0�y<�ca�h�RF��TJ"�I����d��86���	�n7���)#0����w^�*^Պ���d
�@?]����j<3M���1��Y?hҙ�u_�+zj�Hֽ��˫�J�G�b���1����*�l���00�v�đhN���H6$��#_"����YhR��2D/�?s͹A4�D�V�t1 Ň�V�M_����/���o��JR�n����%d�@����ĵ�&X�����x�ɺ�2=%x� ?�<�����������Q/�b�0�8��3�v�7�b��'U ��m���4緰���*9|CX�����f��Psg��}���B�q�0�	`��j9
�ө���wf�T�`H��%�p��3�>�DUc�ME;x�ͻ<<�Std)]���mkBwV�)�J@��B�x���c�j|6��P��2���?�'_��>����s*���gD[���$�/&��F�$b����v�`�5��✆6D���%�<9��Љ�5�5�XlN��s�8;e�� 3E��ez�i�'b��d�=��5����R������8�'y�6����j��=Ru+��P�>�IR'�61�+�3�ǃ�ߥi�n#�y��嵺H�+�SS�u�	:!�A\�����s A�̕�v �|�\K�_�����`��0

�^V��4��9�����h���'(���ǜ�]�|��m��B������~/V�������.o򒖷�|&)�Z��yX��Y
�/��y��C��5��)��QJd?�Ή�����P��Rȩ1�Ʊy��A-��9P$��D��ށ��|Py�q׹JW��u�T��pE߲tV��,	� ���k���N��>�c�wW:vz��fh�V1�'
tX��ؔ]MՍ�6iK�+\1c��f�"�A��%
��
\�8)�r��NK�V�3���ۘ��e�P}z�du�Pg&:��G�Q��;�F��$L���B��5o������2�-�@#U���w���޵N��4�$R ��ޓA"��R;�0���h`�'vR���C��Y0?.dQz���Ak�,��a�r^� l��oC�/\Y���:D�ˊTG\��(�*OEJ��ܹǬ��tcIb���f�c�.��Z�o��bQIy��òD 4�)L�p;4�rfȜT�]={{�~w�s ����2Gv�53�o���#qe���Gŵ=��T�cҼB� ��̝�?^y�Y5��wn5-���e&�٧3`m�H������i�5�l���x�-	0���wN,t��*:��O�`�?�ϝ~��fp%�~wɥ-C���� ��9Ѭ�$����~f�,M��
�4���H`W.�!�1��|�EpD;��S��(�#��8����
p|�D�d��}��q�� O�uA<nT��Gy�cL�-
�)�K!�-B��;�C��38h��?Ż{�u2��n&��n���$%�#/�95�\��o��ߩ�p��ȋ�i̿̽���삥(�)����hˑ�f���JFm�]_���~E� ����� �����RΚ�c"��S8��v���jk@��e��i����	��Ἑ2�	7q���c�M�buz���)�������׳,/�b��<+K��p4�Q�K	%;oqX��y����#:Q��=�i�3u�~Y����~�-(^Ç	4�A���7?b5�"sfa�Bx�I�M#I�P)��ɂ��h�p�&��G�Q��kv´��A5�����3@�/K��Y�����^�?]У>�����Aď�h��;��iGO��(�*�&@�\��O���I<;_����P?��O���b��^��S��r�m(�Cu�y��ʉ<��"v=�3���K��7�l������E��V�y���@��H���8�؝��7�]���/�4{���$Mk��|�@,�M��}mh���vP��+��^�(@��AuE���0`��KA��+Am�`�Ks�b}�Au&k�F����|�ɬ%�9|1;Y~�uGZ�	 3_�L����QN�3�L$*�=�g�Z�����
NR��~���f�g���{x��ù�-Yv�%IU3Vhgh7��r����� ���z�Q���R�&��Ӭ֊"�֐l��o򞴷JyP�c�^4�c�*�{9�<7BX�HZ���Y��j;�Eή�����te��2Q�g�G��b�r=
|/��b�C�"6;�,[�x�&�	����`j�5�4,En�eE���S�v�
�-S�T�#I� ��@�ˀIɀdw>��;�d�hAk$9I�<��������h+�ᑹD�YQ����4�P�J��^�ظ��ɞ���["���*Ű{d� �KZHP���mo�Z�y��<�E����V�>��#�V;� �FE�uC("��g��L��A �2�b���eH�+ăX�Q�L�Gz�qT"�cή���V0�/}�8��)���v��.��M/]��=�r5�"9h��V�Wu.��@�Ǚ����5���j����C�����Bg-��4˹<��EƝ��G��ؘ7����Tй�i���X�aǜ�T_X(�0r-�7$�6��l)�Q ˡ`R��d��ai���9���qK� [枓�ȱ$rg�6=1<�;J���i�[���D��S��>8�XK�/�͓����_~�S��AW�C��:`�w�WE��)q<��٫��"#�d�J��,��M9m�f��j�f�&Q��p�&C��o���F�2V�%�?�tR+��jr�s]06��w�PW�z"1_Ug���)�sQ��C<�1V����Ѵ���~�F��V�AN��wV�,�4��8�˔v��I�c�Þ���A���n�q�+�'b���&����5έ`��ӛ�j�4���z�i0�����8�s<�*}�dz¾{�x��ԯ�q��\��h�S 4S��1T+x��
+�0�n��>oI�J%���{W�l3/
V���~��B@o>���%̗Q�/[�O��C;U�NP��荿a�Y�����hQ��ƪ�H|w!����W5;���r��ְ� �g��_q:�Y�W�=��4�d�ܤF,�I���Dͨ��Z���ꄍA^@�y��d�f����|3�H8<�T�%�9U�`�N\
{�j�H6�`�q;�rw�VV<�,�5h���H�<�D<�C��T[w�SL;���yS��]؍�!��>ol����Ǩ��ɚj��*ޱr��8��s�8cL�=�hR��0�bW�	���J�N*��߯��m]y��N�+F��ː���9�h��h()ٜ.��>q����n�{p�BsS	_����U��%�����5����
�}�H��Х�����
���+�6.�0y�U2��-7h ��Đխ�=SAN�#y�6uy�a+�j�4���Ch-Z�n���B�ɼ'��&�-�p:��pND���(���FY���`�G_ՑL� ��F��[�wۻ��}�"c���v��܄�C��]�G�֊ţ�06&O�CCZu�A���'��-�ExгX�g��ں�')Ѓ�mpk��<�4�n+̒���C�4�@ߧ���-���)%̳�]�F�B� *��?����Ue�v N��Z��O�����A�
��:z܁)̊�^�j�(cXR�N}��o�+�q�;y�F�e=;L� �GDzվm�Hz�Ճ6a�TĒ��� �qq���j/�a����Y�񯳆�ƊQ&"�v�Z�E\�Y�m^asA�8��XC�'"?���2��G��y7t��)�rc'3��	�;1Əg���U�k6o�(1�&F	���1 �2��AM�}N`�7�*�ן�����I]�n]�B>�u9ꍝB�$��%�9�	STl$h ��B�~-�mt�����Lu�[��JLA����p����xn��'�ë
��ZJ��I���j��Y�p�
v��3�mmH�/�� TF�f�	��ⴳ3b��@��[�����͂��=�P ���|�����U ���G��`iam����.n�#���|�!k�&Λ���I�}�Z�m�2S/�d���ֽ1Q��{
=����r�� gTU�.�?F)���YNi�l��u�����\;��to�	c �+�Ǖ��̮���V1@�G!�������3�v�:Wp�tC��Ըc�0t.���L�m�WK|�Q���̕^�Eg�!�y�a��s��ZR]��LdA��/i�k�b��!~]&\�IpD�z�=3�Ҳז�P����� �vmj� �&�⎾��u2�C��pޫ�Zu׎OhuIot~y��QAp�7�	.H�p0�^����q1��U�-�ו!��,^��R1�*:��c+�z)�d��u��&"6��F)#/��:qPA��b��C@A�� u!�U?�4�6q���@�Q�S21.��i��pr%��h/@�Q�'�:� _��џ@������A�o� �]ۈ�`b��V�c9�.�gF�D%�����9D��x�v("��yzY{Glݢ�>����
;DT[rAV����=+"q��SiX��p9J��Y�B�6^�s�5�t�&��u�1gm��'(�l2�%;�b��H����d����i���}��jMIY���/a3�k��ІD~{?)�=�"T��x�a�)��a.QcD�5+��:��[�����
�dm�f��Hq3q��.����[��.�D�[%߲%�?{�^�/�jaa��󨰯�m��J���=���S��a�W8܊I��j��´p^ٹ"F{vO�����*��� =Q��~'Q��|3ϿӰ�� h^o ��z	��3�kf k��l��`޺�-����]�0��cj�\k�����Ս0D�3�R3��H�y��'��M�<�����WI�Q�\�?���,%���Ux�`p��Q/��|?J$�<G�*K�M�& X(�������魤�ŖM^��+���=�-�1�~�� �,=��*2��ů�����Z�A%\��ov�;Z+��@��Ao���Vt��$�o���D��*�D5Fjކ����K. -�3����f���p�y��.��!i�6�爮Z(BY���p�!nF�?�����L� 3�)k���H�qYy���#�A3��U��(�#�������n��{!��u'��`l O>����m�	\#��|	��$}�@���xO�5M�[�͍���:FĀ�i��I�[k�1h�~��ܡ�^��G�Ka�װ2hߚ��y���:@:�q����	O&2y�н͹�="�T�U����j$f�Зu��bc��89��yrՕy�S�Ul���E)q��F	@�	��x�j��ŵ5S;ޔZ5z��/./�-R~��+P�%��ծ��S^}��y���������	�"�-@������ ��4sƔ�o) 	�J���<������5"&+o��q�1�a�貿���[�"�X�?��]בâ�O�9����(���0��`��*�i["Y5�D�'̶���E��lPS�$��*�@q���յ9lF@���t�љ�Jnq�˔�AG{��:<���q -T^°�<Nv�#��rk���D�������˦]��c4枲]{��ؙ׭�ARx�V�hz���Z5���N#�gV����p>�3T�֯�U�����H��~�k��ճ+��%DH�V�r����L�YHG8O+�"�	;���6�%���<3R���{�q��MW2HK�9w�c�z��,���C�n�0�y��w�Z��?H�=�%"�t�۩����C[��Şe2�� �%�r&;!���H�a"�4�֞j�Uy�őkm�hLɋ��hQ�?�;�Mg�io���ux��c�G�#�^N`J�����L�
j��x���>٦�#�h2��%���3�9�B�f*H�s�:p�ϿAp�{�*����^���T�[�d�Bt��A���L�N�Yd���^�'��p>T�KU�a���l��Wu��UN!�x��G&.��JCꁀ)�@�ɓ�����`}���BS(<M5��D����{ՠ���k�LN(A\5�ӓ43z���<2;YYz���EA���t�0Q)ݘ�	��#7}�磼�X�I3	]�s��a�D�z\��W%�AS�������z0�O�ߣ'�PΪ_�:N���"�C�Z`h,o�;���_^A#�������~�Dx࢖�/�%nݲ����'�x����z�iź���!��8jZ��\B>�{�c�(���&� �����ѱJ�=�J.�J�𜻳k���KI�铏饮��ف�|XU�h̴:=^$��9AU��v�^ET�i�L�lr"p��uxM��;��艉�q�sU��X�F���A�ƽh/Qߞf�����ff�}�T��ǃ��ި�����H	i�>Q�� H:{ph�'�ܓ ����9�4�Q(�˟�^���Ve2;�
���8����j��F�m�j����i��U��H����
zn.}�
�+�w��Cv��bީ���s�I�=�U� �z��t�n$	d��n�^�k[�o>q:K�k�5T[���*qt���qd{�S����C�(8����O���l�Z5S�`�[W3>��yP�·�$��Ҹ,�` ����6�a��1�ߌ�ȎW#h��qH�{�L۰�r2q�CDk�^e�vCE���H��Ag�(�"�}8hK��`I@ &c5rv� h�r�;�i���m!=O�Hz��U��Ob[w���|�D꘮�,Ȏ�7>�;WO�*�?�!����71�UƸXtK�y%l�W���Z�7��������u
4Ӱ�O9s��^���!��W18v�g��_LE����C���)+'��yC�®��0	Gn�r�&��	���\�F�qe��B2�JȪ��*���( 5Ù`�~`��>�F5�$s) |^���uZ���G������7�:�7��ņ�pߏx�M>��"EٙIN��uw�R0]�.&�l�������K�"ܑq�}�v� \x��7�V�>.�9�_{;�ƽ�q��.�>��t;Zb���Z0��H���I�ߍ>�o�/��Ǵ��=ޓ�-��l럠��@�$�##�E�#o���F�r�!2����ǖܶ��Ȝ�,Q����wէ�� 3J�e�y�{��J�i�_�7^1���-� �T<�ff�6
1EI�#��4G�ݦ���=<� �+YN����]�3���*[��d�1g8&�,�GR�h(��']E���`R�ϏHfx?Fᗸ-B�C�"�]g���ֿ�;[l��a������N�~��T^dF�v6p���_@.�H��
k�j�Ì�	+��,�Ι��l�+q�żez�;�
3n���y&��l�V��]��J ��&��
�^m��aA�}wa�Dơ�wx@�yQvWok�gO�7"��?R7a�+E`��)#C�;���"P��6V��i��-�ζ�h\�����e�k�Ƴ�X��2�B�d������G���MR�{�?�YU"���/�:�,(�pB����rX}.���#�u�/{�p�>7�Ɗ�����^=^�!��Q�E\uV��^ј���>�H�\:��F����@i����J�j���p��$;� 7� Qd؂�$�`��߾�/B��7�=�g��2%�5�d/
l�[?����ft���!rd��Ͻ�T�~6��Z�	d����pF0����WȻH�G�<�a���㤝g����OK�����f"�(�nR:����œ5Yx_�f�pT!�?H{�EH�A{~��A��e%������=�ޘ�O[�i����s$)3u������Nɕ��Yd�Gz �V������.I�7�d�Lf�uL����w,�X�'ֽk��˟p=4����.)�Ա�E&�?l�p@;Q{*����$q������Q�4�Q5�ּA��	 en�Q��󂹢`	c��d?�R��YfZ��b�B������������w'1��c��٭���nO,w�b$굣��}�|$��.���E�t���u���1��EF[ğB����=)K	�Y&CU�_��a�P�EAF��I�9]U�(e'�H�/���=��Š�}��S]�iT�¡���N�b6���V.��R�;��X�}��(Kj8� ��p�D��a�nw�p����a#_�
W�g}�,���Ox���2ھ�[�m���s� �)~'T��8:!� �}�U��Q�_+�XW�GDh�0��*9�:�l���O��;t^�E�2�r�d�}�f��g�m�$�O���e�~�ʎo*�>���"6�{v� ��j�������Q����Y=���Ї6TBb:,| �0�Η�B66IL^�$G9][%�����J�����!w�'V�mW���}��4�܉�K���gO��U �����o�?���\[�o���~��
��������̐�:�����詼�ܸ��$:����^�
]0�l��L궻��K�)�oG*#�ԁ�u�������'�R�S_����XjES�X����������3�]���Z�X�UѶt#�������/�d���Hs�\K\c�6z�p����7[��
�J��DuZ�-y.��h�˓`���kQC؇ ʑ'��++)�Xs
�'���cC<p�O'�'5���%���!��}J�[����Y��fg���s�Ի�QK����E%��|j�ɖ��e�_q�Ŵ���J)$)0�i�,4J`K�f��Z�\�T�I�lBt�-��6���� �����0�[o�@���`�;4�w"Q?"9Kݗ����:)YiX�9��0L�T{�fYg��{�a$pl��l߷1I��-3�>�G�Pk�`��Q}�:>��<-S� ��j3�0	'v`���)�ݨP��S��-�"t�i����P.��S�Өx��eh��7����W/H��ZIJJȇ�-{1�ڳ���y�p�C����@0���u���qE��0dןw�m	�X,�XkI4g��L[���e
ľ����E�W�
2Wb
��7d����ǀ�P�ҴbWUF�=؊�#�?V�3�6���i���i՞�����Q����6�<HP�{e������z4'�C�e���{�@�g	��k���q<�DS�U��ǎB�{�p͟�ɘ�ҟ ٪C˯.�_�������#pj�28��c�^�+���B���6�
6����@�/�J�-��'GWZ<J��K���>+��Kd{�M����B��·Z5A�M@"�ϔ`Z#jo�Q8܉���lm�ruY��Z.&�7�/>
~oȊ�I�-.ŝV+��<��J�H��79�N�1
"�zħ���g���睝nBy��lw�31,;,D:��@����v��Zi[���Bͅ%מc����y$�>U��z����Ջ��1!k����xm�s\�ar�*�&��d�����X.@4i�5��`�s��y_���~v4�,���9ց��1Ao؛�݄��W�fV������)��#���7q�^�4z%N�!����Ë��@�`���$��`�AZ�����F�y xU�
}�����FB�<��Y�J���*�I����Y��8|h���M�����򄼋�.^2A�qSh����+�0mL 	�߯�މs�c+�dDϟ�Ĭ֒�{="��r*��h�!�G�jzO�����)4>m�*ij�i7 �ד}�Ҡ��8Eo�l`�0fP����s{jh#�;-ֶ��VXs�t#�:Ԡ�_=��tB��6rl�?�$?�S�]!@Z���\��؋�1��I�\���f�0Y��ܯ�(�C���%�%;t��) �Lh�s�	�)�L�tEƫ7�)�IlǪ���ј�ݸd��4��h���#��#�-��R���XF���/��QV�~��}t,���ק����ki~Nx�Kf:�/'�v��fN1�[�_�eF�쀥Y���֗Im�(��v��RĄ`�.���:��Yܵma�d2}e�(�@��ވ��J X<9m%Ɇ$���d�y���;�g�S��|����֓��%����7�$��ڝ?$�C㳕b9��M�[���Rb�� ސ2ꗙT�Qܷd۱����g��ŵu)��'�LƷ&a'5��U$�	ji�jq$�E�/��u���2���jjF��O��"�����mr;u��4��c�C�����ɴ?5����~�O�����2C�������H_�*Hr���i�K�������},Q?�|�gS����9?��a� �؎ՕKw.�Du��U��̴�1��P��#KQV�O��Jw��Fv� �;���h\%�1-�^���"*MNΑp%�qя��	��"��K/�ᡍ��L/�!I����X�@ �
*��A��d�ڹ2I?|ȵ�dF���+H��ޖ�_�RG!�Pe����hU��|Q� �Z�d|�J���̈́�mF��qd] ���&�i��8�%�\��ܭ�ȕ���n��d��~�8�'uѥĚ�vp��jW)��k<��-/m�;���Xz�A���fRW�ɼ�-LaÆ�ӈ�*o�1�T��oT��A���e�hj��D.W>�0��v�}V���)��p�Pp�B�?�˄�5���C �Nב�E��ʠ�����H�O�4XNv����b�������>I65y��N���s�1�-Ƃ�"�K����$��@�ډ��Z^�K�s�LΊ�4�ƨ��r����O�1905�����-���"�6{B��h��3������x��~M�i7��k�XP�l�	���,x���gF����P0]';�
�"*���%�Aiy�R��G&�2�/��#�����[o+���O7�1�_�q���UWd�ī�c 8?����nV ���� �x�|�r�z�j��S�|Z~ p��j$��oabeD��mR����kƊ�!C�W�ڤ����xәi�D@��Y=?ԫ�C�B����,�9�դyA��������r��021�M�8�����5��
����2��bZ��m?+�����w��'7��P�*�Q��<������W����SLf�I�=}���f���Y�~o�N	�c��JA����BT0���;��z֌n�J����0�����6+�I�?`3\�bz�О���}ҵq�f�D��'��7���6��/��p͞h/�`�8dw��CW(�( ���
7���k�-@
<Blj�0(4.)w�RDݧӗ:/o�d�L���^{U��h�J�̓�yN��Y���N�}��ٵތ�e隋�܀�{�eJ���Z,w���W���G�}�`������rP��GZ�,[M�>F��0,Ӭ�%E�g�����rӽ O���OgqQP�҅�_����E�ByN=K)�"4yć"9��������GjF[I������f��nm	�C+����66���!��1#��>�]�~�2���g)���@��C3��sT���e��+���[��s��kη%0qac�j��@׵�-L��]���T���^Ƚi�ٱL���7
�Q����ϠM�n:GYr^,�aP�$1�$�|��Б���)��V5�_�ts)�����%�grZ:�#s*�%�xu4u�be��|�*��a�[?�*A�LW�p����:�-�:t:�񼅉\h����F�!L������Eԓ)�cJ���d��=0d'IK<X��;j��t*����K��� =�!D��M]�����*�_�*]��V��G�f:�����O�o�牧L_@۳4��=+��?f~@��[b�4o9� b�N�R��s���0�؏�y1
��D>��X*߶"���5��(,e�x����<y���J
#¤f��d�	Z�����tI|O=M�D����:�$���0�f���O����J4`�Z����¦cQkv:�<EC������gX�����-�4蜼B��'{\�!oF=�%����ӧ��M��=}v�G9T��Q8�bO<P��.ʐ�&q��A��K��ME�&H>�gi�8�ݱKB�9�໹S��IP�\%fb $}���N�6鱭��)n�y�j�nÔ�[�]|�S�+�˚�J���,o@<��k�=�K��1O_K~2�]���"����0��\u��������}�db/�$�m¹��-B2�f롆����x�INt�ڲ7�yj����,-+�u���,�H���RZ�rm]�#bΚK��o?|k�˥�w ����%��tԺ��"{�x�-��U����:2}��:�:�V�r�T�JIO|?;o"* ��ۥ���B�1%�z�++臘>eSޑ��S��
�g�ĭӉ�T9��OI呹��3������b���W���\R:��5 ���K�I�]o�ϹG���%'XȎ��nX��A#�~ʼ`��)pI�V�0���2�0��/��^v~A��z^΄�jݭ�Gh7�L�p���zX����B��lVq|��y�ֺ&������Y�qr�:���zA��kߊ^Ϧ��mG!� n��3��a���JI?�Q��Օ��fu���YXrG��#SՃ���s�(I���ck�+	� ����dW�V�8��ʴ�m��T��WP8�Ęr��n��	�4�%�AL��̩�P�NI
k`�����4Ao;�C��h��o�v��P���B�%�s��Β�$Q_ׄ�!<t�sZ!m"�U��I^�[�v�O����{�DNb^�X��>��
	#fL����:�3o1�����O��]$~��N���B�Q�=Rw���C�f���M�@��uxp+:b�]��z��c�#,���w�*�V�{S���%��,٬�c=���w�o8��0��g��[f�}�X�0���r*�Q�w:�=��u/21��zvJ��P-��ڶi���E����^`���%���.x��*VFe�U���7]F�t�\����Y���#�7;�W�n�)ɹ�p���@���/bGX���'���1sn�nu�]5Pɶ��TB�����ٕ<��+�Ɲp���-�nT ��u��R�,�F`�P�Q���})ێ"���K����ح�QP�}%��b���$��ZO��!��x�j�����)qAz{K��B�^�_���k��&5���hy��u�+��}���@^`�cta+� :W��w1d��]��I/�^6�!� p�岫�M�U��X��o����hv*Lċ�ۅ�LY��-H�ɾ����h����?ʈ��m`�b�6�6R��n����`e&E�汐iL�g�:�O�f���i��Q�/5膓H�2-��L^?�_�PQ���O�U��h6~�PxZ�����ތA�Jb��"E�s�,�J�P�^��^����Nm�R�	s4	�:y���u2�j��^0�S�	�����]o���3��'�s���.�r�ה�a_��/T2�� T�E�Kv�MlKPqDX�����%
Zo��`���"�r�yy�h�n�`fP�WL�I�G?�k�����6?	�%Lo�t���w5���[H�l�ƻ}-�	A�!���0��S�j�E��p��8�LP\������"�Jc�Tb�]�h/�vUiZ5)^�3�i���T�b����?����P�'��}�1�t)��R�x�{���Z�~��uN��y4
�M)n�v�e�
���(sW��3ѫ:���uaFK��Q�c�`J���FA�ʇJ���=�} �}��6�\����_�� >{����4q����N�5&���X01��D����}���C�ÏDK��/��M���Y�_��-�b�c�]�J���m��^�J�d#�?��ϭ�����e�:����di�����{y�ي�'ٗ��I�Ռ5��Xj�Fj��t��*i�.hYi'̃�ic'F�#DI)}�浭=#�O�yL�AL��+�k�U��"�Ekǣ�EI*z�]�R�ݯ�J2�'�Hr����Ū�dB�Or�mG����9�w��rtVsF�=��@�ٽO$oy�$��Niw �G���ݟc���d������yx,����D�։E�V��;p�X��9̶������W�(�����'��_9�G�h��g4��u�ž���;�Wo����+����޻���Gۛ�u�T;-�g���k����j@�v��Uq�g��A��#CZ���(��3��w���1�=jF�oMɖH(km%�1ܤ�ͯ��[�4 �p	�k0G��)h�x*p�IF����M6`��Q���h}[RA�8h�?�^wĄ��H(�3i�2����coRFmT/��|�p���A�ըj�I23��>4�sj���9V=�{��<k$Ҧ����ZX9Z�,���g@`o�	���I�*BJ�1:?Q]��A���TBm%�ו,v�_)���$�����W��}x�I/���v^�ܙi+�6�������A�o���B���u��5@[7N]BĖ,�Zf�T�l/�27,�n��<�	��4|a�?b���{_�!9�w�_j٩�<��a��Z�7Eسz�X5�	��o�-���ȜiKg����>��`G ��J�G�#��O�~1�h�e�`b�M��޺V�t}���ןxY�U�	�D��ވ,~V�2���]br�BE����AI�%�� ���t���v�M``��!�z@[���h<j�	�8TL�ڴ�(���,�@v�-�p�E���u�����Y�<�Ѷp0+i�g_�Y���̧hZ��^���|rZ7)b@���;Yף�+q����F�Fԣ�.���z��.��"``r�b��%!x��Ӄ��8��ܪla�m�V]�nG�JR���`���d��l�*�C�Nr�{�����P�fF�o?��[���4換-�����%��nR�5/�mUЊ���J��j	oV�4��̓�y��C�b��*jbH%�ߧ ���U��B��"\L�s�j4�x���b &�E
�ؗ=[�p�y����v��OM��J��q~kR��,�Fx�=�	����J#�R�L>����{]�C�G�e-{���MĄ6��{��Qז�I};�s54�y�_���x��BH��;�ИI~�w�3���醴)A��$�Rp��:Kt(�4��9?hwKO}�em.7K=C�J��h8�����x��V0�`�lZ�y=|N�Cx�����$hG`cbr_��	��#ɤ?�Ydo�`=C�n��@�	A���h*�W8j��q�E�cP�I�e������'���<�$��]*ۑn�
Y! �\P47t�t�ab���o�<Ӷ�tl�,������3�,���}p��+�A8Up�̲�.ô�^���Xg�#˖�(��H�T��iV����)m^5�:XA�I� ^C�X� �b�0>�s(!$A�0��|�c�d��J7f=T]Ä^�H;��|8���5�W�5C����f�o��	�uC��X���\˕Âm�.�`�i���Z9 �P�rI$��OV3��kJ�m�����{��NC����1��޿T$��n��.��L�nC����eM���k��4�����0-pnq��3�@�s�a��Ֆ��7�;A �������X��]�L`�>�%Rs�p1�kz��w�¨֦E�]x>��I��>eCE��O�B�ҩ��e�R�}Ht�-�T�1�8���ך�g�M��-6���E}��´�Vr�k��˝��5y��m�dS��/��|J)��t&"���;�h&)��i`{���
�[��M+���0S�B���Dֿ I6��9���>���ReL�]!Gs� 2ڼc/��]nI�,�ۇY�������=����� �m�6��!>��<�
7�q��J�<����"7р��y�����n�e-��_w��w�-EVM˪�=���g>�׷̀�0�`���G�BL�?x�9J<Ȅ�XY�Ӯ��H`>���/�w�g���`��6�ē�x���@�1�[���뻩Tڃ{��p�w�-��.ȥrGHq/�!,�����:|���7�N��qL�˃��	oz��#�v3�������k�ل��a4�U{���5?�+D�2*�p=9@u:�;p�v��`92�@^��R���D^��~E^��9'w�tCt�U�L���#Ԑ�X���$s�8�"a���X2��z^���G���:��h����t��� 욤Q��|], �ʒ5�P"�,D�!^��GG��d,�s>�j���'	W�~y���Tri�$�5����e�<����1��]� ];�N��Ci%��H� .��=�^_�T4 <cw�6�x����f1gb�؇2d��SP��W�J{��{7TF���n ���8�۬�L�:��#@+�p�2�n\^P���)���?��Q���{4?v�l�GA�0[�͵�����(fH�ag�^攦�@K.&�h���IS�Y@�Z��_63�xHn�\oh�vIo�δ��˂V��YO'B�Jx9��]_ ���w �L.6�jxyZQkN(���5��[�+Ѡ����ǀU�1OL�rK�~)� [����-)H>��7�A!���o���1��*$�<_w-'b������U�h�Q3����_<�]��ر{>��o��<�7��d�/^�5��nZ繙�T'5��51�ۥRğ�1�0���Dˣ���x/���t�#W���V���*t�J��^/�:o-�ca�)q�4	H�ȽJH7��JknB9�B�AK,��(�i�C�!"{ 9��:��#��1�> N�-�RႦΕtd��YA ᵳ��5`?�ɥ�8}V�zLQ���ȼ��YOm�����*�_�_K\,Cל����[�v_���ŧl��e�Ab�M14��h�ww�c�|7=�g��(���F��_� +{���Yq�T֓�����䪚�U��7�7��|w�:�o� �ظϝj�;]=^���sN���2~�-
f���WبG�C"�H�c��{�[�3R�<m�+�M�C�pFd0����o�'8S+`����-���P&��l��,�a�u!$s�O��n�O�_y��j�Fiє_�U��\��"ZЉ�7Y�g���Ѩ�1�X(%Mr�7ŏ�K�q�9o�H<�Zx� ׂ�hZ5�T�Artџ,��aA^��� ���l�IA��>�6�8!@��+�R�k�_>%չ�|��P�F����>KyWN�J5KlQ�9���X�jΦ������ĭ�[�lf�N��ݣ�R��\���qR=����Oj�&�v��0ǮZ?��g��9{��+Z�ڴ�恰��{���"��9ˢ)�a��]�<]�F�[��&�J48��^�:� Y�`�bʲG�w�Nw�5t�j!ZsJpJ<���wvj�;�yʇ���MC��4�GWyD��?�.#�Z�xc�v�<�K�Q��z�8h���Ԙ����3b��&rR^JwU�a�R�"Ӱ�]nʷ*Ǽ�#�*'�I�OUV�Zf���|�]�ԛj�Xyy�^f�6>b�Sp&IO��&(ݓ`r2��uMk��C%��{7�����c�?��U��r/^���\::�<9�?���N�G q���Vh��WkM�ݞ�ĕ-x�u��l��}$k���+��U���l�����m���"dGqk��t�歪�k�]�^ߥ�p��];�� = ���*��>�?�M������x�Ց���FƊ��������{�̸:�?n��7�pBi�'գ.7�E 7�P�2B���jIT�\=�VS|���X�sZpʢt���c�����q�Xh{2����,��������4��K�eMμ�B	�Vbt� C������U7K�)fJ)�FS�KF.�ԃ$�. �e����㪄b���y�u�(E �H��Лe��c캁���+�Cyd1í�h'cL��P8�Ī�P���-F%N �%!�4�����ͼ�GepH�2SI��ko��m���٬���m��z��3t)�'�f��2�I�}]y��|�H\�&nL�\�vꨌ�F�j[��7���%�h�X��S:W|�k�b}	wz��r�C�M�\CI��eK�=�p�l;�� ��:X��' _��ÛM�E�"�����x�+P�1�J��%,#�60�B]� ?��S71����ej5�H/؂P9��m�GK�6�t��VvM"!��;g�rQ���J7����Re�ը�sJ_��ܪ�(�-��S�]�S���YzP,�x8�l{a�J�kP���,p��9:AO�R������g������Ir�浪�+�Ja�8(���{,�֔BEr����M�V���������k�	�����00��&T��7H����֊S�����3/B���x5A<A��k�t��^�AP����Z�$-^+��U_��3�aL�&��q� <4��3�@�Z/��Q|��U�����6K�
�Ǯ�����ȅ���ە��8����e��#�L��"�����~��ͮ5�r�L\Wh �T�Z�#�6u}�<��9�$�+,J����� ��V�FьV�M+���٘����y��g[_�嵎�j���*�����P&Wh Ü���6̏�Tg�]2� �1@a�O|��@G��8��*���`����F�j����� ��vOw���Fve���HW��>�&q��B����[�{�^�!��D��	�R�A"?�n����8ƎQa7�R�۞�D�g����T�8�]YIi�-�~�d�9�%\ ��$�qm���{���D�uױb���'~�̑/�ZcIS;g�����7K��$x�oa�p�8���#����B��rr����5@z�T�'��Z�����+�+�v�.�>�(z��$�"[�S���i����.��B��n��w������jj߽�&�#8x��S��f���eƊu�Zv�I� �]���y�5��Ȉ�����ȃ�<_�;q��<�h@��%H.QL/-�'��o���'��A\Z�� g�5uSɄAS��4w"�kfo�M�*�<��D�xv˟��T��Tn����|F�{D~B��P�G&&���_�La�P�_U�E���#��s�1ʫ;{^��&���=��� �B����KJ� j>%NLQD�\3*�9�c�f�L�g�T�V���z��d�����	�hّnh�>��g����n	�&�J�V'z��������R�>��D����O�{�F	A��:!��_�:2
J��C�ܜA9@
���jCo��6�٢j����ί�l, ���w��:�5�"��|��%������lZ�l�Q�`�ya���J�&>թ���Zw��!�C���T}ѻ�U~�a=��a�=m��N��a�n�bx�uw($��Ȉ)�]F� �דk �-�}:t>�#/=m��שc�V_�������A��Н�[�R��&���+{�$Z	����������W����tu�S�1��YX�h�}՘؅�ҹ���0���wB�o�7ChbDR^����.#3i�����:�S>��o���
�ݳ�%kPHa�kfAcwާ��Rd	
ܥsi%0����Wtv�?�C�@�? v�=-�Ǣ����-�ն�H���:��_k��r'�m�.;���1��4d��˯�c�I
��v���vIj�y��� �%�ҹ���-�{2�`Q���U�Ă�z�P�t��#�pԦ����0�g��ti�����V���
��զ-��׈��l1oC�r�&	�^�a�z��/~�=�-;d��0�*B�#|�7��k1
�������,�z$��p����B1��b8!�C3��ݶ�|V-�	��Ҧ������Ь}�nBy��).�q��Ŕ`���$����<�Ӹ󚶏�-���"Z�J��L�/JLy�?�X2�U���2g�,�ZOa���?܈Yu5r�����V�21���,��0�Rl����ݶ��S!�28�!�i�&���a���*)�O1�n��/�N0*����f�+�5x�
Wm6�Cu���)-��*?�� �/2���!t����D��Ȑ3�w߾��.���x��A8W��n[��)"^�iM����Ux��T���z�S���)M̉�SP�i��}���+�J*�Z���P��h��ԃ�u�'_1L� ���e3��1�{��i�)9��nA1��C*�*���e�0���D�Gֆ��e�����j[�'���qIf%z�iΌ����`N���2�XItiv̾Ķ�i�m'���!�B_�^zI�/��;����vE�,��l(�D��Ɵy��n��e�$�,4��V��Wlu�
�(�����+�0U�rb�ahJՎ�Mgqp�]����%1�zk�M-e��"�xo�1X��\k�"?y5��KE��Cy�芌�g"�w%�%�I���
W�t�-L������d��s��W@��p6͹� �e�<.��(D�{�x����)_t"���_	Lg^-m�V�ZG�IB�K�|��`+&�R�Q�q$s#7H�cv���s�7�<o�E�"ve��&/��`�C`�D��},mZȍ�M�=<|�*VS��44�ƭ1�o�T�@h;�97*u��R�/�O����Gg�'�&N�y�F�wxk ��Mc�J;hg�Q�/@'�W'\�ʃ~��_Zr��T�f�ST�*�L>�ז��p��zl릲�= ����Kx`rO6��"]Lp�xi#]���m� P[�J���~��JD��^7�7�����9�Uܣ�����c�֠"��Z`AF�"����kH�x�hĦ\�|����.�ǐ�q�Kld�fq����n��~*b�1r9E�})f0���r��/Fs��p�'�Lk�B���c)�Z�5�Wn�����О��Ҹò�H��4 ����l�_�ޙ�v�v�&��8&S-#$Q�����C��z}���YH� ��t�ah���bK5".�и���<�S'��v�2dX�uO�n�o��2:�ˆgm�
*��Ti�X�Adb&�R�F���=��nF����f���C�9���kFS�ʰ��������
?��E�.<+@�w2 �ۢ����Q�@&PIn8�C�Z��&��n�pD��{z���j���T�6Y@��Vz��	;G��S��;������~��O��ߧհ)���_�����UFI�O�w�p.F@��`r��A^�f7_b:�*��r����hS\a��E`@��g���M���=�x]�P�ɤC.כnO� �!F������f%�d����!TY,�Ey\�����2�x�0K������0��A�3ɓ��h�S��f���i�t��>ϘH�-
���n0B�	��|�۫��֐�:���O����(�rV�swd�!��n�<!�
AD
�L"�=0��| Q��~���I-3��8$keoL=$�F�Cq�>����A_������MmUX������@������AL�	�<}O����צ�*�\�Gt��F^P�oe�l�k����h�XA8Ӿ;�Q<�KI�AGM�R��ܛ�s1:]�t�Q����	D�=q�N�3J�G�g�����y�� ��Q�4H�k����aiL�����-(Snh�>yo�i����%5�/e�u}ɣ�C�.�0[��LڼG\U�C������?iY�9�K���&)�]�)2ha��<�G7�n;�aC<&�)�U�dH��b��1�Fq��' ȳħ��hv�7��q�1>��Wz�U���Sk�Ԙx�W�@N���¤�w�?0��d�9}e �ш����i�tT��G��R;l=/S����\Ϝ�y@yN�!.P�*Ԙ�o�@ ���V9�B(��{��_JR�n�J�6e�n����u�*��i��y�X�¸���M����72�6呥�#[v΃H!p�yd��0�x��v)Xz8�.%H�)j�Q/�
wJs��A�-�3��fۅD?��yT��pYtG0��ʦF�J!񤧹,�C\�L�>Ϫ��G����/�]r{��������=��B�tHQ9)�9F"� �Q�ðU��MY�
��ܔi��dj�1
S¤@��<���2��=P�/;'�J����}EL�voЭ_{�E�c�c��$ᠽ>P2ɫE���3�'�s�M�y�_v��!��w�ÿ3C(�� Aȁ�~��x��s>�3�t�r ���߳����-�놨���������;F-=�����[��uU�E�f�.P�|�U�[@\�a�q=�Y�4��,L95��3Q&V�@z8j_/��~����0�(�!��ZsM�y_���}I��&ʮZ�Ԏ��nOAD>5�\��!�&��\+�o��%���0Ϲ�xQI1ɓ�&=�c�a�� ��۵`n�0�PXYC�I.	O>b��иx�Y`n�'ӻ{E��/�5�=����@��d�\o�Ԑ�pt�ز�F�`�9*�ԓ�!�{ة��^F�&�Ȗ�z��$�aǧzs�2>�0Z��{�u�Ͱ��i<�A�m��a4���cP2�و��ys��*�~�~�ΊɎ9�M���8/�tj�;CSǧ��09�u�#�=c}�47��ޘW<w�I�O�����sr�䏭Q��t𨁀#�}}�&��3��)�S�Q���3)�8����)c
�5�"���G�
a����j_WHlQ&���p��LL���z�&t}Zz�Q������|b<�);��L[B��)K�Kl�͢�o��-�5��(e3y��\S� a-x0���a�pDgh�c'-r��ԊH%�^>z_t�
ȱ���œ[�Wr��Y����4���� ��������M5�_��&�� �*'��t]�e}���RK��2pY�E��.�6~$g�\�MIIЍR�M*�vA�r�o'���������oI�I\�9��h|T,��7�@�'j�C�*���>u��*Py6
�l�Iq�JmN�������bz|b�w��5+�(זl�v�!ɹ�=1L8��m·=�˗�{Qnhbr���8`�xƖ�m&@���\ ]m
�@�Ȕ�,�fR��B#J}�G8[�)ſ{��-��4��߽P@zqMl�C��0�\?j�D2�YL,J�CAŸ� j���B'�O]$K�H��E���I�Y�p�Z��c��� P�@u�f��	��<�Gz*2�I���;0)�$��t�k�w���S!�w�T�~!�Ｓ,��Tq��%7$\<�!��ͮ�8̪��|n��^��e/'֦	�nc����@�d1�� ��q��*��|��7�v��!-˥��?��ixk������ʠoz��7
Z�y�ۄQ��`�y �����Q-���������D��C������,v0�9���S6�8��_N��G�����[���G�6�m_�5������'Ыp�\g�"���V�YZ�`�TJ4(�ZpN��2��?��
݁e���0[쿩m�?�c�g�NO8<pc>�"��tY<&�U�k�y���E��8��0�0���:-<���6���Y�n/?�J-���[�[A��� �^��6&v�j������t:������ax��>�������Xx��7Z*m�L�4ҀsX�m<���O��R
$I�H
�v�!@5^pB�Z��AxL~<Y�H9�k_׭�cBB�g�� ��|n��pKx-$�<T�w��-xb���┩�|���Rp��V��T�57��[���ہ{��y*`}"��!�2 1�� Y��5��0�����v6w'0F���� ��1�9����8�d4c�2���מ<Rʘ*�r�U{zb��r<�p�8h$�}=S��7Pyꩠ�Z����f���E��1,.�J����)���臐)@���!��"�@�||����6�E!%�<�
� �aH�ch���(7�SPY�pM�T�K[r�bgt׭t@���B[ͣ�:�\Y�҅���dsMJq����t��̊��y��M���A�ڣ���l���ahoAm\F8����V9�����Lh%���,�b\q�Ql(	!�(kC��4A̬��7�L"�,�䷷'�����e��H�n���9:�W�3�s9�%p��[v��/�'i�:ɉea~�g&�cc��_���_�#*V�`��ֹ�g����v�e�7�ێt�$$d3#�:\W�[R�H��d�Ƿ5"r܊G#4�s��۷1+T�߯jM�����e�p�i�ij���b8�/�rOE>W ��'2S���-�|Q��nH��r�Ρ<����W���grHV�e~��Lk�0a&�'�ț�Sq�IK��8���k�.�|D����O3G[�,q�|��s��@}���S�z%��@
��t��%G� #��O��q�yt�me��<��>l�:K�u��F+.��F�(w�]����/�#��
5��u.�����F�U���ւ#�bg�Z�ó�Ψ�01Ǚs}[O}`�2��"�|���6�#��s��ٜftvW*�QSN�4]Ӑ���G>87"��HV���녘b�pf�Υ:ɹ�5�Ǒ�B�d��Z�����yf�l6∖<�+�u���$o�Q�WT�*�����"����ݿCno������$��]؝���4_Z�p��%��A�e�� �]P-.�^�������rc��xy�
���1f��qј�P,FGHq
��)�vb/�)#K�<Y�Z䴀J̐��Laʷ��m�8I[u%i���oV�E���*9ڙn���X���$; $�~���~�����.B�gt��niIZ�p�(E['K^� �EC~f�����<��ؾ���Ajj�Hynn�."[�6틗�ǉ��DP�Pf/�1�����>F�h�#���p�T�ve+fF��2�m[��E�~-�F����%k��������cbi7�$5��!�6��h��K�[�H֝�ap��ùV�&�v�:[X|"�W�_ͨm�VK�gB�j�,ӝ�E٬���qEr�ކ�4��_�b�n��$�'������hB��p����^5�5���Q�2�9W]	R�ob�8.TRt-i��t�x��yhr'j3����)e�.�(%�رѺ5�漲={u�j�O���Pd��tC2�x�J��ʇ*������8�Z|?]�e��SY��t�0i��U�������O��
��d@�0��ᄜ|�>;��8����B�$ڋA1$'5{�
�١����Ð��oN��l�dD��)SV��ȭ!��K���묍C�{��;����8��/ȏP�b���˃��\IP_�t�^�{�u�XD%a���y������M��0��G\������pBo���P`�:��� z#k���c��d�oS��
��?�g���ڽ:����~�F�f|H��Fm=�l1�e� 5
�W����Ct��[�gtkN�L!�#��Wbb^���I�@[ͳ�N� ^~`4�Fӕ�l���B"����qP\���0�=�}�w6��Th5[:������It�|e�&�����o���\8:���#����?���/�ա��[�t�ԥC��m�S��� sMKX�/YXs��� �PS!L,�x�󀛃*b�����!��gat.fV���PB��k��0=gA����3e�g)�H��u��M55c�FFc�4f�>�JC'�˅C���װ_�v-�r=�s�%,�a]LQٿ�F0URΞ��Lu1� ߩۨD���w-]��`�W˨q������7M���v(��� ������Lx�訝�2��|mA�6p�XП�
�i��S D� ��-{����`���kD�s¢���;�i�K�,�Y����@�ŭ���%z!P0�/��s��?I���b��Fˣ�Y#I U^�����u<��_ B�N������Qӝ���(^O�B7��k3�N�&9��J�v����� ��F�d`6x������?�5�_��c�MI�8q�.��Nq�X�KgD�.2N�6Nf^{�af8��������&,��[˶_骎x����_���r`��C�)�� gw/A�UpW&Ò��>�=и%�|2���5>���O�'��ڬןa�I=m�ؑBh;T�?6�X�D`�/��q⹋����b��Bj���B�]N��gB`xc�]�������K*���܅@�U��(��Zu�92����� � Q=C�+Ɂ�[soEm �5g�l���kP�$��81�j�c>���S 2�B�����@� �0J�Z��Q�P�K�vEs�7�m��'�g��6M¶�6�[mb�e�w~-{�BP�|s	t_mq���n�KLP8���=�=On�����l)�9<z��8>��oT�H�����K��ӎW�B�h�J߇���ЇdҠ�� Q�a���C���.��˟�{}t��7�c0�V���^�a���[�KE�������N���,�f'�lf��'�Y����un}�ߴ�W���
<�i��ӊ`"(���d&s~���[b Q��EE�Xg#�F(j�p�����-絔��JQB�Aկ/�Z�1%����b- uW9�x���!�H�Hv��V��e��,���'S�G;����6�n��Jv�L��X=]�~b�����;L<G��{�P��PM��J0�(Ջ׳�o*hk%U�EV��TJ=��,v,ov�>�D��m�L�,چK�������q�e��X�>c%����t 
Qq��X���S��$�j��>���E��㉢�۹�O�\�`F��'�k���j&��]���B\�ٝ�]ry�R����8���`�����$Nn!>f7��#Vض߻w�ЁR,�Ѩ�(��V"�Hίg]�#��)©oK���{����`�E��FÖ=�ϩ^�I�I��WG
:��8���f�G={0
�j�]V��<%qx^f�Z��~j%;٠#�F��1s��c$��Z}Do�V��~�([�Vj���/�NH��0a�V����#/�d�ipo�(Ѩ҂�����V��bFOH��":�(,��L6j�'/�i[��Gb����s��4��ɖ�WO�}��ʅߋ�I�Fz#���	��#�y#�W��ry�P��|F�֗z�>�ݺG���"���7���û	e9dK���	��^8�]oӈ?��
d)p���X��*U1ә�mF{��|&���G�M��~r�)'cWr�:|Ui��'h|b�"G$�Y#�9u�!l��������J�Y ��1�/�h#���i�qL��
O��M&��h�]�;2�0�G��#$�]o�!�^5��/4�P�AS�Ĩ�ְ��u���:�긢�j��Y��>�h�s�!����W�z�:2��T�Jq��^la�^6�.YW��9S���R�8�&�¼Tg����=�'pH��;{�#��	���,�j���f���}�)���ó42��~D^�L{�7�t
zτ�5�w��Wt�R�����[��!�6q���
y�9,�v#B�����]ar�`��̏-���N�X]U	��:���H'0��$�k�����9BG ������`_!�/<�E���a�y���C��L>ëi�����q���y��$�)Y�Zљ�e���*_(��«�f�ea��^F��!��`��>:{�s9g��͆�f%���?J\4�xd���G�Qv�Wr��h)��P������\�C-%Ë���}%�Ǆ6��y��A�����˛�N�ީ�.9uޥV(� ���M�]Lл[�#"YN�)~3���
ׁ)&�<�������ı��n:8���Ixg#n��C.)��SM�~����sn���|��D@FU�C�(;WG�a��A)�ACZ���A�J�te��㿢�<2�� �\��`�����V��y|5��I�Cl�Hc�z�5��H�ii/��=�һ���Y�����1�Lx�3CV?�V4�~�|h��ϸ<��9��Q"�\�$��z?U7�����<W6��l�`pc��G�d��?J�if�
[�,&g-�xu��!K�Gl(�њ|��	�d(�ڭ��6�gE�St%�f҈��G��.8����}yp��0}|1�����Oºz-�~ˍ�A�#N
��]����/���P�]a*�c����Ys,P����Ev)�3L��j��ōD{�ןնU���W{V�H$K���9�9QUU�G'��Χjh�R[^|g���!��:&�X����&�v��%1w a ]}e�8�
5�^5��|�Z5�-�����D��p�5B̧"ߴf�Qw���ؖ�Έ�!P�v���#2r�I�F�@=�u	}x���!����1��O��	a(�/��j�4O��v6�Kio�>�g�" e���y�~�����������7��|��B��{�a� ��ұ�t�����$D��;��L+7$�l�S�79r<C[u� UG��=!������K��MH�]���4{Gr�����N�0��.Y�h��c|�3�Jm����;�^����8̸b�VƊ[�
�r��J��q�A��:�B��^�_�j���qG8c����]~�zS �r ���A�>�GD��[��%����3�?��H�C�Y��	ǝ�6��n�Jj�����d�vƖYq�$o��к�%��E�f�v�T��'�[�x0�/��^}o׾j��=�����~b�q�����E�ߍ?ӎ۳�����9�T�cc*Xi5���PRh�0���2Oo�^�b�>�\&����r�8H����խ2���Hh����_���"
ih��>���C�e�g���n��H���t0�YR#���*���Bw�߮�џ(���r��G�slr��`~�$��6J���v�
�1�~�ώg��g��+���Ei�ϛ~�/E�����j������M�=V���\3�꺑p0��k�n�f�L���`��	����TE����aˏ���v͘G@���&���=�Z!�]��R4��mfu�m�F}A��#ґR�|��� ΰ�BlR���H�ڬ�%Nd��`��|����,��("���`~�-7���5���L �g=�C`��˱�2@\�+Ĝc	�H��~���Q�|k���S��1��K����i��>���+5(���ʘ ?�џ��9�g���}ɥ�������/XӢ��?��t�����R��-�1(
_�Xn�����O}35`sʢbr�)ZOM����%�e~���6���H��e��`��C��J�||���"Z���O�j���
,���<�6�tP�~�,��z��W��4��3�b��8)7g�ɲ9R�Of
usKo��Mɡ�c]�ф>9��u��]tv�Y9XUS�G���L���ܟm�Z�h�@EE�D�&ʩ�E�z�̛}V���mI��^vuw��A�ᨕb�A6b�/�Ɩ"~�U���7�kJUR"��bH`j3�R_ҿ��XV\{g���ݗ����hO+����3]��l�ެ��0|�$a�8�C&������GhM�V�1�����8��a%��ݗ��)�7{)K�0Dd2z���je��b.���E���Y���QW=��Or<�*yp0!�\X�d㟓���>P)u}���q��ǣ˚V[J�Y��9���c��آ�(�[њ�=�r�b;���ҸDT|��U@�Q+�����4e<����8}�'H���є7�G�=^��&h,�&5���1ÕZ��Q�N���={j�֧��E�ԁ��)~o'kM�����x��Ȅ�7�3;��~�G�6���Ր�@xU��{mӥC�sK�ʖ�\�c.@�Ӎo_r85�!e`�h28<�p�X^�,6b�h�6��l��_{�)��܈��N|��Mf����B)�O�~7 p�m}�������� ���������U�M~r�VL���XS_�Y*�����=�m|t��5 �>˪*l������ C\�Fvk��!��AoyɡYdf������'�b�g&���%�Jd(U�e`�+�>� ��KJNfN�c;�<֩�O&E��۹ⓖ�O�vr�8�U�T*mA���N�zˑ�g�gA�I��6I���8����N�8�Sl��2���R�R�J��.�e���a��ᜡ.k�|wd��.��Gh�P�e5�3:Q�������컈fX]%4�lv� ${�vNZ!̻^��Ehf������?	_-)Yj�1E�-���Q���l�n)�������W�QJyN��a�g���a 3Vcr�.�	�����,I��^�^�� 4��[p���u�?0@�_�/�a�Hؽ`�銡`����n���zt~D�$
�v�a��-!#o�wn� Qn�t�����H��r�e���`rRӐ�J�������H���f�.=Ig�}̝��w)�:��F�O��N๻�]�F��G�7.��55�r���\R�[����K%��^;�h��莮��̎W �e�p��p��㭸�Oֺ�Ϗ)p]w@����QN[��%u����!Q�������>)&mB�Z:�v	5���8��W�+�=��gOJ���pZ5�Y[�t��VY�b�l�%�ى�j&�|�A�a�=o���\N&^%���K��v��)?^�t�N�b�P��dWw#��V/T�+��
����}w4��%}@i�3{(���Ȼ��j�:���4���X�-�!䖌J�ı�P	@�ǁL"bA�iy=T��L�Ϩ�����Z�x����sV�V�,�����a�/���	�� I���g�Tt5��2�*�b|�ld�O�/��^0���MQ�5���E<�x�S�I�����*���k��r0��t���	,�B!H{`
�YM�GR9��4�7k�����T���� �硓����.P�����A�_���x�|��d�%��T\}�ϼ�jF"����\��C&94yo��
��("�l�%�O�:���vcX�Kh]]ەZ��E �� @���L��z
3�m�L_�o��G�zY��6��j#2=�D���p��h�H�^ץ���N�5�w[�f/�� �Ja@Ψ�H݅2{�:�}���^Dn&��c�T}���)��Y�8Z�T��ـ�CFTy4�K�5P�hM�"�l��J��=�4�,	+�_^� ���%��"�I�XGs�2�M��o�������~��j�����D�������������-��=�C�W�I'�ط��+�}Lz����e�L�ԡB+��D^QQ�ܖ
�t��#�䠛�,q���y�qo�A�iGI�h,ǵ'���S��r���T��`3�3qĂ��U+���~�2���Q|����a:(i���^�-�Jw'ˏ"@v�{�����|�d�^m�ඖB}��	3��8N�PZ��d��S���]\�eM T
��=�TEd�$�ew	����j�jg�.q��1{�[m�
�%��M9�1Z�ȉ��£��j�8�d>a�Ā<��Ny3�������Л�����q���7�0nBK.D0�RP���S�Q@���b�N~��h^TWO��)p|T)��$�q�ߔ F��ΊM[��+���m�Ѿ"zҨj��XF���̮"t)�,ѓ����b����"�/f����*D
S�^˄#�q�z�+�K^��"�M��Q�}hׄ�p������. �se�1�i�����v�.�Ñ����j��xr���FwA]:3�́�G= ��2�q�p.���-�k��Dh,���^��q����!�3�ݠZ�a��f�hY�*���j�+��S_�N��z�.Y�ܡ^�`YE���HyE����99@}�$�;2韟	OyP��mW?�f��yr�Ŧ��8��1곚�לVf%�˔���Uտ�F)�ަ.��ׄ$���y��y)�E��7�8i�%���|�$���Q6O��f������ǚ��<�r-�
�yȓ �!u$ Z������@ܰ����ty3��o�e cT� ���}�$�G:�6Z^�W`���U��M�5�R�φ!�����a�u8)�W��Q[7T�N�~��am�u��s<e�b�+Ùsu;���u�r^f�)��wv;d���8��Չ��+���A�M�Mqr˲�/�":��Vh�6��1a%����S�eF�#Eyσĉ �m�v?g�.�1��܇}�j�`5/�᾽�&f�B!����Gz�r���J�.DQ���u_k�$��0|g�p��A��LpUO�XW�e��
��=@06���ԭ�@a@����t�8��A���Y�:��� �fTk?^�4[$6b��nK�h��,�AF�Lo�&(�C蓅��q6�{�?�����t��9���7����ڳ�+X�!j$��Sf��.k�pQwr͡\G��7�f�$�	m�;Ї�/8A{�aG�������n�y�`�0��7���c�ִy�j��Ju�ܐ��[	�67�&"�EFQ��#Vm������i�Ymܻ��
d�)}du'�J�]�e�ic��MCluL���O�P`�@�.�:��Q��ە? ��:��T�ͽ�������B
��2N�==���Dk��mmު������\���;��ϵ%���H�#]�^��:Q���Na��pnW+��5e���q�#F?1��]��րL�|C$�����=_vW�%L!�����luwE�X�1�싰��+$|���ֳ��rq
�=���{�(=̝W����ZrHr�p�. $/�GY���7.y�U�(�Y,���1����$[r��,�M�փ������Div�yY�� 4�hs��X"~��M�M)��p�_F�M�h�X/�-�RҜ�E���%�OU��6R�XZ��O�-�8��<P��by�x�İ��#�Gw�v���uFѠt��[7����?b}�c&׀ft�,��UeNT���P�a�|'x)��:כT����n�B�Q+\���E���y���tsG6�q���,����q_��*��d��"��qMצ>�̔?p�0D��3�(�5�u��������ӊʎ�ې�>�=�"*�`UN�G?@�<OזL,]ǓS��[v�2�ި!M��)g�������a6�Ïl�	_�w[������Sh������q���c�.h~�N�[X�:'�P�R�`Ɗ_��肑}>9��^Jp��g]��(&5�dv�9��-0���[0��MU�#6��3�C�ϐ˅%se�_�G��t�ς	\ '����-�`}�ҽ���pB�q_�L����2�v뇲[<!n����b�E4�sR����}��?�n�Έ��!AEr����֊.\z�=���el�&w)\j�ޝ"�~(!����Y�l�R�F&�N��SPg�0{p������l^H���Z�ciN���i�u���>C�7l���y���8T��*%�?�k"�V�m"�@��_�� � l����=�i�@�ӟƬm ���Ж�͕f8��W�ę�����Z�j�`���5�|��ԕ�9����k<p$�E�A1�&������&�I��C���wU��l4�ݲ�<�1(��P�	�~�W�d~w���u�7�c��ϕ�5dBz��s�Y.+B8�zB'�W ���U'�����°��Ԃ|<�?�M���B�0���W�7�(.�\���F:\Z��ȕ0��C��?Xwb]ai]�б�c�
8��Cx�,�eѰ�L��!��][s���4�s���i]�t۰E�J����}'Q5�A��Ί-S6/��t�U��ë���}l���8F̄0&�R�߭:���[l�Ѡ{�P��k@�`�l�'��?,��V;�8SY���$��B�+�Qy�g��.Y�On��4`������c��׸��;�X/����E-�R�3ć�*�:�|?�~pTr���{�/�gc�`�g�-����`��7R8 ���E�n�*�ĞƆE�jY����L��^�����(����~KZ���=���sցc�ɗ�cCth	�~�_?��m�-��j�OB͆�WJd)@��*\#�t�c%NC��EԿ{"�>HUkI&�Ow�z�y�Q���X�� O]�6j�ƒTM�"��{�g�1����g�x�<�˂�8�U1̦���]^KZ�3fxվ���h%m0��x�YV&bKTD�[��6��Y��/%y��{`s��e�l�Щ�a��zc��+����Őw�=�E�'���ne��aw���x��6��p��P���z��~6�瘚O��'_�m0��UmX�mˮ,��.�_V)��=��t����z�I:�z�//`�[�/�-v6���d^<�Z�#�>�ע�{�߃���rCa#�?��Wf��#OGY������ �;�É Xj��Q��RUv��^��Mr�|�![�h�٭�ΰ]I�CQ	]X�2�I N�F��
3�
�!��ې��i(�BM��"�(�,D�k_��J�:���5}}<m�-G��%����k;L�z��q���$�9�ʌS7�V����������c9��(���|�(*yO��̚�"ѻ���(��*�iTԌG�4�qǮ7��� s�����Z���ڋ.'�
4EcS[���qr��A��:���h����K�&�L�=E&��3��&�y;�]�S��	&�Y]6#��	� x~�����8w1��iXE�ƓDzk�N�EM�.�0�wrU �04�t�K[��aE1ͻ�l���?��*�Ʌ�6%��K![��y�m��˲tv\{t�P�k\��30�=�ȿ�K��^f��|��D^}�{��'txZ%F�0��J��p�*a-
ҁɶ�=3���G��ƕ"��w�
����j�5H4��sJ�h�*-ǫ�`��-.t��0jE�p77W99dl��_�6�0�q,@�i�jݐS�B.,��z�bl�*�b�ݬ0[��:Z���N.F���f��>f�+�E�DJ'	��	������k��>����_������P~<��2��Ŝ#X~A0��DC�g 6�`�c�`�>���������Q�E�[۝�!�`U뿂C���q`��{C-�P�z��<	1�J�x\��f�M��a^�b��K�d��jn
�{��[��=4�'߾6N��8��!t�?�;�3p�@�ɰ�tz��,l�X����А��Ћd����t�;�����[�CE��xOҌ�4�8��"ezt$�Kqk}q�\f��)�<����S��kHr�=��#{9���m���m�!����MH�#�N@��DڹgC��� �Y���؏��S���q2c��"�Uy�FP��ul�kR��Β�2��嵤z�����Y�|X<�Fy��
�I�������;:�-I݃~P�`c�L�1���U�k��Ju�~���pѼ/y��)����1�<����~��v�>�5yJ���8)��nٻ�*���O�����9�I/���O��VjaV��l�k�w*����K�I��Gp2!��Q��Ɨ���i� J���f�
�,�#�\�!1��Z�gk��ɑ��BI����&�]$*�H՗���6�r���vQ�����栔ʜg�������u�IJW.ɽ�`�B�e
���"[3�C��<f�[�Mۍ�R��R�.��6YI~}1����}�,�f�k�l��+��!��\���|���7󲢆2���F��\,͐`r-����D���Gp�h������3�D��
	&��Ўg��;�Ųѓ�K�G�.v
q���n"�/M��fKԱ�q�	^��]�
��+Q��?�9���cћ�;�e�N�g�	��m�;O��%�,K�\��.z�g������Lo�A���A�K_C%D�!{z��=.�lD��VS~C�I�����  ��n}��y�Ňw�&�W�t�'�p���	P�`R0�уK����ݯ����D��������!]v�{x��_o)����ʙ)�/	%�g�[�����\���t�f��z�M^�,�������n�����o��L�'�>�w��(Ƭr,L���G!�R��y��	�71q�l}9.Q`�%D!�Ɏ7ϧ<��v��28�"U�-؆��h���ݹ�K2����ݫ!��]'dQ#��	�df�)�svX�t��!���>�{'�J����p��0�eМsK��g]���L$�J�<�e h�:Lƭ
�oİ�a�z�߾d���.bO�4�P���j�P�I�{��,t�L��i�5��Qw�A�2ZƠ���E�����c�>\�<ᎂ�2J��[pS��1�P�}|���t�r�Ep��\�+>#ti���ah{���s���Mp�������^��nL���F��6"6��©j&c@�4�F�T�+W��Ec�vPu�$�=�*��e5�H��J}�:�{q�O��n�֛�>�s�0��F�Q���KΘ<qF��.K�4�f6����adPU6��Cږ}a��L���Λ�Ҥ����K~*Ldr!T�k�a�����c�I%��om�v��6l�+2�|
Y������m�'�
�������=cD�K��Ӟ��c�B�Z���Ks��<`ľϏ.�UG^�q�j��:IlM�t�B�yFAA�+܌�G�a���:0ʈhdb��Q!���L%+�/����B�Pj��`������"a��~��<����M���p���f��<V1���=��B7�AW�h���z��K������<��g�OX���=��㯾&�!���� t�d�ޑ�-�IR��Bmx�0y��@(�*d�L�5mҿ��hݲ�q�d@�R��n\�������Uf��`���3��<���]�YU�2B�$
���������dH��K����˝K�X�,��i��R�E���ݞL�������j�x���Ұ}�KaG��W��G�mzX��#�?��_�[+;sq�d��[ד{I�3��̛	�S�&�=M���S!��vs���vVہ$g��Y�
aU��1��h2��ݨdq|���7 ��]Lk���_l9&41�h�lޛ�^Q�ۿC}���M�j�9����%[��,�Ԯr5�͆Q˾�-��g}�� |�:��t�ϑd�W��]߮�֯�> <�N�P��XZ���|~洒Y��,ɡ��J�W��~��f�������g�c��+v��ܯ�I��D���%k׭^��|���%�DK����8��7)�t��":0���L�y/��GXHdp���"�v��Q���ϗQ�G�W04���b/#7\` Ji �5`�z3�7� ��m�
9ok�x�H������0���\E�?�f�y)��y=W�Y�e
��S�7��Bo�ZVR�5&p��n٥<-/W��ࢊ�L9��^n��� H�Q�9�k�U�Q+�{q�v�ry	yA������(�1լ�i!r��e#T�V�^;iH�G<l�i��!Vq�qݟ]|6���|�=����qXm����?��ELRX��aeB�p��s��D6ׁ�f?g��t�|m-� PXب��P�b«pGr����Y�:�� |����6a��������r���U��Ԧ�����s�B3�� f��w@rDbIOy���&Sv�qE�z�;S�PN��*�~n��ݧ�<��6��_KT�Ў�=�"��|9��%`��Gd+엘v	J��5�O���{��o-^�5)�_�LN͆U")�PzH�����P	�U��s��k^�a>�bE|�N�#ЗGMX�.��WE�fP�F*�]5��֌��"WH�-�[����˘�*�Y0�'����?�����ޗ�R��I��ف����x�����#��c��+�S�7T�f�DJ9rJ�nO�k����ݧ"��c�zQ�bm�l[G�Y�����:�`K�)��r�e/�wE�j�����fx{UU���S�wrZ.�^P���>��*tn���o#Y���j�7�x,63C7m� D��1
;[.K�/��\4�8�Z�'�b�[�k����vM��	>eѡ{d��@��%��
^�Ɏ�~"%7Ȼ�U���9��	�W���\��L�R�)���"#'�-�KR�Nͤ�e1�����Uy0�����PK:�.��Njb���_�jL�@�S|V�E�'��wl.�#0�g��'B^b\ePxK������A/;_�=�R�Fq�I�<{�:���P�N4I��y�^����*�̕��殗����=ØW�{4ظ��c�o��^:jI?\����)�9�L�?K��Aj���0�����C��t͍��G����R�:HS�K٠�밎�-�7�֚b!�B/@�5<���J	C�/�T����i�}�~)�3s5a�G#���V�W�h��w��$���L�?�7��PU����\��xˢ��v_Ҟ�k��GԀ8Ph!��KufN�P����H9l<t�	N��g@}��fp�SƬ�$r��j�]������=*{�����ͻn���U#�PxhnS��~Y��|�j���>�A?K/�L�!�_��?͢�~�v�0�Ki���戧��'�4֏,v-�����mۨ�8M��O"e�Sg^�u���Έw*0*�ld�옞�Λ���~��/K_��t�A����}��PH���a~��4d���6�WW0���%������G�j7#X��� ����g�> ���5���mm�5CD����.Oltj��h�|�ߡ����̕��6���_Q`��-��Cl�٘��5l�q$��+;{�1=l
��.&G�/e�	c�U"�q?v��7F	�L�_�������sw�ݏ��A's��׶�g)֬��Թ�����G��?���<B��:A�C�jdv�Z�>,&z�T��(�"m(^�e�XqTese<]��D�6�tboe?,.��1�NU����^&�����Rl)��ȃl沱�g�������U F�L�~d礄��Od�*
�eo�k�ְ���u/�����^Ez��I���S�E�`Q>;��7<]�#��8�������4�D�T}�
�����h~�~�v�3�|����a�U<��Pם���)\3��τ�,v�}t�y���i�h�#��3H=ͼ�����o�֥�	�����S���������B��f�ҁYY��q�v�ж�����+��$˴1]�����T>�v{�h�	�4��,R��4a���#k��W_-���-YSW������q�L/���:|���P��{�tAjk`qn<��в�;,M��d�tܶo�O���W�Y�w��><N��l�h~^�	����4���AhA�H��j�BbE�䖛��O����S2���^>.s�F�C��A��`����6�?�|����F�c�H��D��v�|ESr�ei�@m�z�mZ��@yӞ����!�e /�vߥ����_ʨ�\=���AXb�G���yI#����juA�"�����L��;!QVy��c�X&%���[֮��NQI��N�kX~e^�@M��a/�앭fּ���?�"6&h�j]�[�y�p;�^>�V`�9�<*�Ob� ��!b+���D�8�Pׂ1�2�_Bo�y��^���w!�YN-��JՔ ߶hŒe��s3"���q�0�hjM5-f��R.��0?�Q�),�[�/�����R���~����ݚ�=�T/�N��1N��,咿Ɇn(Q!:�TS�T�r���e�4�f5492�E�gT���z(�0��C�S/S�
=16��ӑ=��?J�� �%Ƹi��C�biom���ͱ&�/.ܾ�4�[B���
�E6�pD�
�CZ7�1F�A�Y~%i
_,:�̛��IrJ�G��8&�܇>p��I\�4��1��#2���H�tV�(~C����g�k����~:�fgk��M �sf�1��A`�B��k��W��M�i�{=���5\��5:�)r��s���պ[UF�0�m�u��YX��mٍ
�����J�+�ci�T�|a7-�?�A �:Z�^�HTĀ�S�R%t ���iеç5�p��zwx��umr�1�Os$��#�mV�ӔT�]��~cdQ� ��$%4Kp���L����c������9~��)�N�A@��KX)+7�߄���w{����'F2���7���Ӳ̹ף�`�X��*H��TR�?�����9�h�}�+�T��1̅�r�5����|�����ޚ��]��l<"q�;�4���H�5h��H\��ʠ��O��}w�����4`'u�sH(�'�DlE��?2=��h���s�VEA�0�N�!}\�E�ra>�. 3Z>&��7&�Pz<��F�H�-m7���+�j�M:Y�B I�~�z���IՎj)f3�o�t�w��z�hrc`aX��A2t��?|ۛ��������<�k����J�YO���f���.�����'|���]�>�ϿKw�3�z�_����o�����/<���Y�%S��8��R�q�_�k���yR�p���n,�1I����L�<P�gb�.����eYt��x[�t[6��h˿� ����Z���_��r��ִ���E��"G��'IR|�����.~��f�P�.���/�i3��j��`�Y���֜{G�(��R�L���m���m��'l�.���V>��p�Y+��6?<�����)�O���q��T�󈄚)s��#jl�ަ�-��e+3a��E�4ƶZ}�LԊ0��V{G��;�RU`j;���t�����gR�]B���sp�@v�"���	�뽰���i,�vD>��sʤ��N0JQns&���Ֆy�|������]�;��?�y��u�t=��F�� s�6� �1q�AU)�������!��uE[?�`=>�Ʀ	�&t�q�ҹ5�[�b��&?ޠx��`qٹ4�o���X�硞�#����M���n̋��A��\�b�C�!�u'��ܨ�m�:2 ���Z�EZ�h5�D�9tށm�9�`H�
���aƟn�`�B#�b�Q�)*�	��6��e����2,�K�C~���&%��0^z��B�y/���b���r��G{nY�KD�c�E2�@�ln�_ѷض���yi}G��6�'�r�7�6Ǭg{T��TE4�0�,��ʉ�9N?��(e�#*U58?��}y����F���?��I`[R�mUJdג��i~-�\^~[o$Q�9_n��wn�X�����7�u�Բ�ŧI����:��!�?$�*���f!+�6fۺ&�ǅ_�6��F��#����F����U��JE�:�8� �E�)�����4�;"�ohD?b�vܩ��kq�(���ip`�M��92�Qϧ��욕s��8}���qh����ބ�E ;Ǝ�����=����Xm0�7ԟK���F@�G��,�a��]̘s1�>��p�#�+��^��X`ASi�f�N��s!�0�(��g/�����^� H��|2D�;�oW=ht~�b����Y�Y��6�:5�z�|{�4Ye��Ӹ��y� H �uU��Q^J���Ss@���	aJ>�4���uMe�ؚ� g����;��[#�N��c\�.|O6F�kݖ<�Ds��^��e�Q}����;oXh�(r`��yQξyi�D5�&�I%0����%�&��8$-C��뾺�H֟�"3�P�v�$�8P���9��18��EW �3�T�ĢC(���Bħ��yN�Ty�O'G>��d]�:U�^O�-���}_���5wJo��i�:&�Yk0����*A�߹S=@Q�r�$	@1��+nQ6�����(SW���q^F�vj��ф)��E��w��D#�L��.����:C�xR�k��ڔ��fW�N$����� r�����#�ωϟ�sn�X�Vl��_=A)�ͦ�����a��Z�;@p����ov]HC}���"��ljkL���o��pO���}	vĔ����8ʈ�?�WӰ�_��p,V���"r�����gj���P(�Y�Q��5�^b#�$ouo�����$�Ün�/�N�8l�UV�`y� ��h*̰�q
U�X�¥�.�����O��sB~,��LB#y��Q��-C_�&�+]ь#�
L��3�\��slV����^�y�cAL��KK���������5zXd̰�}8��D[�C��J�K��-@Q���-�A���[D0wa.�:�)Uώ�L��g���2+LH����=�+�",N���J܊�o�.y!ߺ�R�xm�fo�\�Pn��^��?/%a��$LF��ݸ�+S��Qq�����iCl$��������7����C�v���i���yiY�����=�<�rO��*FC��#�?~W�y`��/au���]�7�6C��i�qG�yz
����eϮ��Z	_��@2�_�ԍz
��?�lb�J�|������3)�����l�F�œ�������x��TE����;�?�I=4Njx�ػ�Ꜭ�S����qȍ��e���z�ȋE3��e��k<;���|��/�c��VSܔL^w@��y�m?^v�����n����oӿ��H���� @��	+gv �̷7���]��+��
�_T�g���Ǳ�eR ��WlvKB�U��S��=V|�3�s���b�XA��]�ֵ��]�me�v%|@�ǣ+� ���UB&on>�.ZG�L	��ʮ�ȭk�cy�{|�
�ɟ�7���``��_)wa��y�G%8�A��fT�`�{��)}�,�bN �l��8ˁ �B���η�xO�l��"��>��Ìr�HH ����R }s�'OX�7ڢ�`�#;E;>A��C�)��[l/��۶��",��'���hDs�r��j-�c*�$�GaP�D$�w�u�;g����<����dT&BH�\�ἔ�T��!�ٗ�����g�T�6ׁ)�H��]J�}��4%'5 ڬR�Wb�l�{3N���*aT�p���Ӑ��ǜ��)U���G��d�1��,QMA��$S̘q�j�f���J{f�1�RM�.�K<���/f��>��o���H�@RB>jX0�&�˗Q���y��	$5������F�x0|%8�Ӑ����/lb�xv�V[����<<�lK�NaLsV'e�&�:�Q�nY�+�d���]��0��]\�^HʚSm����I��h����m��7����$�u�� /��u���|(��t�zewn�ߓX,<��aS��
��z�u�	$�=���8�/�� ,��^W&�嬤���	g@�����9�0|�����Ȑ䨮�%�:/�l���;#��$��|�5s���7����@��&}�z�$�zx.ь��a��P����̶qFE0pp�t'�jGӍ������@Nb� n�O6��K_��b����ߥ��D��A�����3rXz�T�4H��1ß�K:�Ubş~�{�]���K���!�C�k2i�m�8��cJtvδ�קv�������	�]���j�7�/9�>��f��M({Ѕ����x����W���B����K�vcW�So����8|[Oa�V�[��S�2��(���~����Ǹ�SǊ_N�G弎Jh�C�/)`=�7�K�7C�aLl~����zn�[b��~��ߒ� ȤH���Č�'�#Y��\�os�u�gV�=3��n}Ma�.�wcZ|O*GC��C�MS�K�⫴"Pq?��+؄�W��� �����<��^)�1LCo���9�y3��S\D�(N*k�tD<�^�jD��y�9�S5K��Qƃ|�E"����N�:�yzf�����hE9�jѱ��R��Q�Pf��:��ܘ?�ҋ�;9� 2�����"Ϳ��{�쬊[��>�v�hg[}������o'���q�Cg�������r2X�!�Qo���^b�Z42'<�����ʨ��C�U/����s�����Φ�4���Y�T<��/�Ă�3�@��W�!����u����|���q��jk��Lt�K���7�ѩz��nsN�7�;u[ ��!F��8t]#��n���h�}ż��f�!(�@M.Ə��ְ#b�9�W���i��Ze��	����fѼ��o�e\���#�r��fSX>��|�^q\(����:�����(9ı�C�Ļ���U�cYV�b�U���s���('$|^����,cԸ!�a9����{�0�
�%a�1��(�D�����3�]��L)Sm��K�F���[�ԅ�Ԃ��2�����C�`T.r-ɹ��Ba^�H���?=8�q�g6���6܍�9��;�P\Jy�YGjS��������4v�Ώ�fN��K�3���6��?p.6���1��������ģP)j5W������Wp�lP��r���x��IC�i��E��P�)�Y�u���Mj�r����紆�G0���8`e��BF|���p0��}ZK�v�^5fy�O o.��N��ɤ��a�/�ng������cHsU��te|{�d,��[x�V,+δ|a��\D%��@�e.J��q�G@�+y��.�j�2k��H��r�ʗ���}� |=2�p���af��?��|P����mY� ���	���Tl��lc����{���^(��}񯱪����'Y�<"���s��Z����ȉ3����)N�Mg1��R�������Y�8�l�����N��J�U��
!q�-R����Z�p����C�;�J��(�Hg�d�tk
��2����):qy�SbSHv]��G�gMf��c�Yi���	�4�^�g����=с��La��X^��;k;��>�W��Fi���BLMi}���C�%���u��O�C�Q^T�Ȼ�lU&���_��s�aϊk�K��R�$��g��Y��]��)S\9�G����jp{�̐��Y1�̼����.vNů��PqL߿�?)���aq3۹�c
�8!��h����s�s�.Dn�J��Jǽcm����`�0�%ޟG���������K�β�||Ѕʎ+��
D��hP��jY!�,>2L*y>�8fË���e�K�����]lsЉȦ�Q` �)Cv���P���T'���T׎�*���Q˸�I�B��JG.�j��3��~�.M㓳o�E��%ٽ6�>�Nd}��ff;�k��u�6�ꍅ~QkQT��xq~�����Q����_����D��N�T�j���F+V��A\AvHi�KG�x`O.w�H
\l�NU!��sVX{����L�5��%AE�����yL�ز�Z@�xHW�	�'�O]�?�����V)j�k�Ύ��5ʒ%�%$��b��۽�\cC2~��ʆ�p�t'��J�2o��s�ы8f\�E]�Yj��;��y�w�I'%j8@l�vk��sY�2^Q�,mn�yx�:�o|?Xw���MX>57@|��ۯF�Z�mP<}��).�B�j�P�x?v��A��;��n~��nߍ�n��,��*^YM�*,񑉬`X������W��1����]让n����oH��DLW�I�G�{��]�b�3��ҳ}�=HN�\XjT$'2r�]�|T� �,*NpƠ�}'��>�䬚�틘L����˭�T#t	Jv�nh�zW�����^����/�K'����m�K},*uH�<weЊ����і܎����F<�p�ʚ�\���{ڼ�iM��|�9GE��_.���0(�x�m��Ko���,"�8���),�R���+��l�B&~�=�?X�xx)�+�e�?����A�B�ɬ�!w^�����-���r�T��x ��ͽ�J4���Y0��<����f�w9���uK����*~��}S�/"S�࠳Ο�/�$BA?�W���,���*��.^��� ���g��_i�lnwR,�����Tw6́��.O�ܕ�G#�<�c����Ԧ��5�(E�p�]�|�Hd�`DL�����c��ĩ栺��*���/�!\f;�ҹ�/D ,��XذQ�s7Ls�$�#l˒;���R1_'@^�$k��Z֌��k����+79����7*��G����W�z�$Ձ~���8a`�
����#Ř�w�,Ӧrc�� B����n��ɋ��_ql"�s_�bG���3�R%�l�P�'�$���w0;E�r� �\�NJ��#��@ns�b�A*�ϽfcA�e��ݦ>%jHO�H���/��W:��3�ĪM͎t��}
�%�]#�Ӟ~�a�Nv6$�8@���f�=Z0�5Xu�{�b5A+���н��`���OX�	=�⸊�_��N��-4m�C��N��Qe�KO�GPm-}
�����5	"��=�w��=m�o��=Ҭ��>dC���Ȭb���vg�U�Yްt]��O\q��أ<����M�gI�7�~�2o΅<1���3�{N'3�h�>�'
i;��7�(��/�m���	34��!��a6��� ���x�F&PiW齑�/�WB�������-��1&��X��E�Ρ�3��!��}%73��F���*b\o�|y������ET���铙ʕ�� jK���eQ�f|N�m;�!�������	ZC69�si�C�ṯL�������q��4�RѹD�L�P\�S�����LS�dJ�
��?Q?�*Z����F!���@�vpH�)	�*��IA��&Q%9�1G�S�j�hʒR��r���Mb��v,���ա�q+�}�,�V;�|S^�����eh�:�xJ��R&�~G/��m`���ۅ�Y2(�	�zoPtܨBP�Ho�L	g��~C�Uk,��PV������C��/�{{�l����s,VU.ђ���y�Z�>ZI���o�}n�n�KwA��4�����R�Ii�k��?y��ނ�P/V4Dx��B WKr'풴Bк�g5 �\��m�ޑ�Ч��T�,�����N��	'P�?������:�Q7�.?Pk:	<���T�nO��jJ>�/�z K��\ВR����DS�nߐ��Q,Du��ݫ������\�K����'p��I��8�Q`�R�+���Ӽw���y��^Nz�_�N��؜]}��g����sg$�Y��:4sA����A�f�+@&��0���`q���E*.�Ae<M��|��?|�k�y����*�[u���9������BL���2,6�)4��F~���U4I�p6j$�_��� V=nB�x���^C��Q\���2l�+.�;�-�������&���IO��	�Nn�;�3�^��zqX� �\:=IެO� ��ǋ�F�[���5&���/�U,�종�S���U�\^qI3�:Q�i��v�5=�#�SLG.<��> �"J���D;�5��7Ch.��Q���"�#8�ql���1?��K#�B��� ��ajm3�nɓe�(�:*�ď.��7�ŧ��J��E�1���VP�KԦ^��+D�`���A��
�j�H��$��V��;�[�n�h#A��C���^��騟�Y9�R��S�#��!�ֱ6���R�,�>iQ)i��s�p���A�7e�߫O���[1�  ��ƀL�'���)[Fhh�'�рB�� �l�� ��nR�@=,���"�)��|]���z�-�Ҷ�4�s�y$(iY����d��i�4.+ru�����0����3gɘ�����l��1���"v�_�$p�c4��,3����w46s\M>�-WK�t�P�Ȏ���1Ѕ(g'	�}Ȕ�'T�m֪r��m���nz�G�f���7�tU�����k2$�5u�Hm{vѩ;Q�$0��D9,�DkO1�zf��;���F��=ro�#���];��޼�� �Q�z�;r�?�3]�(�,!K��CӬ��R���Ί��}���a&'e�.�d��Ɓ���'���S���v{�2�� <�4R�%A�͇Z�~6�o�2M̸��O���`��:=�3���(>5}��\b��/���у�U��cA�5���*bTS���LX��t�=���$r�HiӤ�)�|����8��H����ii��Ov�8���u�
8����c����u��Gb5ͤ~8| {vW�]3y:qym�i��
��N�w�+h/3��~`0}L}	�MG����ny��N$�@>�K��y)��J���pHq��xamu@G�$=�����Ǽ���G�]q�U�Z�ɸS�DH�?���3�g�n�صF�4;��L���w�4!5��~���c"�'��;xPW�1tS�!=�;KK�L��kx��+^]l�;�iĴ>��4W�knT��e��I0����R��+%�(��s�n�	�l$ �|�2K�8�)�����M������h�cw�8�I�	�9"��%�g�x*�w|IE����W�A���xav�!%܂�L�\�;2�X)�ĩ5ݼ�I~�e~�������|6g��5��Е㫪��>`ppXJ�7~"nsv�,��w4��c�[��G�.�V1��Z��D3�Nl����N�@~��eŐjh�}��C���+�.<,Է3
��Xӵx�Ր�md�l�ݿ���y�W7��<�a�e����e�ä�1O�5��x���)g���D���w�r�~��c:�8�|����_���U�Nz��mY����S�B8Ŋ�Cf�Mu������ �1���y���,i�; �w�H�~4���d�U*5Σ��و����9l�f'���C�7^���1˵_"r���\�P.ۀVԳ5f�.m-��J��➍W=<�éV�M�9BO���[ ���Ե�{��ZJäʙẨ���S2��\H��}}ͥ�&�fVG��w|~��9q.�`.����Qry+���AҮo��~��e<T�a��y���~�v�g�)�4=:WK�!e�D�qi��RJ]�ݽ�+'�~$�"񟂖UO�wj�&-��>��J�E�MΛҿ�&G�ZX���L�����F
G�g�%�_�1�nrvS<�<�s�a�c�3ף����`��ղ�U[Gi�&��j2Q�D)b\����Um�e�WU�T��M��ʌ�k�� �����|��'@��`�S�jI����-	�~)������.���@;H�����I��@����}H�+���K8B=���=x�JB_qR1���.�j�05\���P0�G:}���y���~��c�F�@���"Y��EI����1/%�!��AŦ��t�5r�2�E��>�圥�K����	�Ab^����;�2V�w��#���}g{�/!����������?_���I�ַrk;!T��5#��xno'T`��s��ʂ2�>G��������}m���GX0y'���b1�ׇZ����>,랖�v��F�1I��L�]����k0��yu�Y�lV��� ���Y�؆vX�f-nи́���'���y���B�/j���ą!|�
��-Ŗ��u�w�B�ټ������&��Eڶz��A�3C��A%�C3��q�!p��p��D}�.���E,�C��~��_0-_��X~�]��O�VT�ȳQ�!�;�7s�H��I��/f�Ѽ.�WA�f]ẀӔ-�)���1�XD<�ds�� j���s�`q��c�ע��MF��Y�x�����#�Q��i�����g����0Gt]=��~F�Gq+L�/s�I����m\v1�~��g���PŒ!A�������d~�C��*�,k�N��z�<��F��Éb��Cl�^��RԿ�i���h�Z?��c-�o O�Wt �3H�,�F*ƅ���g�4����F��gy0i��}I"�8j�	��9����AtK*=c��T²d���_dG����=;8fa��
��GMvM$�v�A�'����i�#8\��C<$Rı�v�'����ɤ�Ru����t1%a~b����4a��Kq���8��;�{`�xf��]洿Mȯ܍P'���R%�6ϴ'I�~i�$["-G�e��$�r>�}b����2��7�q*U��gY!�5����:)ȷ%�]�t��*�/���n������(@��8�-��03�UC�uWxz�&\}g-C�~�9����{h0!)�!{l��TU~V~Wj��{�|K
���,�	�"qt���N��+�W�.�v[b��,��S@}��	.^w��7����!(p�=<�jîͻ��+�O��T
�kB��1�Ž0^�i��s�3�*EL*>S��!�l����}D������hن�y��3��n5G{�s�=�I)F'e�5��^'z�c.d/}����O�]R�����8�����[.u�S�D�� �<o���!ڰ����~�EP,��i��ֆ���~��q��=�?M��^����9d���*�n?ɐ�a��9�����kuk�N	�e�$`MДD��dk�QA�Cfמ���+�; '����2ޢ��+D���zÄ��Ѥƾ=?c�=	B���;�e%����勲�t��=~�����AD��j�a�Α�}y,������Q�e����s�T|É�^T�4v��]��G�k�\� (��w��\�j��2�ׅ�4��-j�5F'O�TZ���NP`<����>����·�c9�\�2�S��ɯ
a�:�6���˲Fr��&%4�wN���I���P�W�`G[!w6XR��
�����U/�!��@�_��y�^s�K�{�v��B_�Е�|,�4�Z��9�6��fU��xcyp�}��Ov8�#+�t:�f�T��p�=���i�=��H�Z<��p��9�4�EceR�`H�f@���o	[ո�Di�|�њ~�0��l�$d��4�� ֓1'�y���|,��?&3p�ec�I'�b���(2_�L�ܰU;�}D�4���'�p�%q�gu��n�AcntV�jaq�d"Mqp*h#���׍��Kd#����X� h5�!,��F�t)M��2���zՈ��ȿڴdwUy�xkYؓ	�Yk�aMh�Yc�5��0;.d��%"��>>�0c#�O�+Y�,�,���j��.��/T��,�L�9��I���vj���?+C�`�TɝII7�Kh�V}zZ�T��F�	�o$��|q[����m�{��\P�ǣ1�t|��ӿdK�Y�����n@�KĤYէ٢6��X�k
41� m���q�:��s�yd}#'iąD��1�)���� �<���w��Ui5̏&v$���3�n<U8@��Eq�ic7��D�l�N�W~���������	%�Ɉ��/@5U	������o���oZk����y�Z��.�k.c���nƔQ��f���@���'��Y���Ae)ǸQ����od��8=��I����۝�W�:�(��h?�mF3ڙ�Z�`XrT�x.̴A2q���z*p7zJ	7��C���x�E-�*HE�~n+H�&�f^i�⨝��2@���h��,���H1��Hv���M��-��c5횘`�]��ﲈ�N�`Eaj���1n(�9���"�w�q?�C�����e;~p�a�׍/���|b�6ǎ��+��Q��cU���VvI5�Է���5"@��R��;*B���y��E��S���#2h�{yD`�T!�`2�vU�8Hy��:Q��iX$�#�ΎV	���ʾ��h�1-Ĭ�q:?�_�эB�y� r i!��X@==���L��+1��]��Ư�g�6.X���R���GDGzQ�P��Ry�b	��}²ɛ�¢a͈��z3q����&�?,��MCF�U(X��N���{8�8�s(ވ�U�r��js���@�-G;�
���{>4���{څoZk���:g�| PY�� E�$�௔�H~�c����O��|=��Y�n^䋪�����A��v�q�s�F5��i'�w
��9n��Ɖ��35&���ɱ ��1VJ�p� G�i�*Lb��DK@�[gF�7$�7r����%�k�X5NF���W����/sH$���h�����}�8����
ھx>���'�^<ɣ� z�o�����ҐR���헠������t�=FRhf�I�� E�ht2,�e_,���ٿa_��@���b���*�r[���f��֛�m��5��{�	WUlh��kd�,��eM����H�M��ǔ����gӹy3i�
֜�gw�X����n��.��?bĈx�{����'����1>+(]f���%�� �*�����m[�Lq*K�#s��Z�㑠�C	�L���m�˚&ʜ�L��1�8���~ݑQ7+vv!��$k�����7>�H�lČ�#m�N����y9Z��l�������Z�|��ۅ�=P5#n���>�ifM"K�?�~��k��y-`���E{��������qq��g��}��͋���-gp`]����m��i����rR$-4���a�Y6�	�qi+����}��qDw��a����˳E0�w�,���#'#��V޿��� �i�4#s�6aFi`��D�cv���C�J^�e�=�@%ʩ����������&��3,z�V���%w�\5�ap"d�:�l���D�F�W��?�A�lY�"������5h��FRd�[��"@Z���u��D_X��O�e
�~�(=6�	�GѪ�gE(&mi[�j�'s���P�/�xu��nO� ���EC��9^�퉓�H�R�
;jYpC��qv@�k�a��ZPInf��^:����Jt��v�m\e�\�S=m(i���|d���z׿����@?��+{T�&ܜ�_`��Ez:݁Z5Z�_.|��?|�xQ���8�3%��5kB��8a�U�ܺ��	<�&.Fi_rmJs��k���b`]X�~������RטD:�>�<�O�����bS�_U0`+GΔ�����nZ����ҬՏ'�rI`$v3	������vE�#����f]���a�R���Ͱ:�`[�L.F��dc��x��֢Ʃ-�]�M�r������j�հ�3�t�.�����S�� c/�`�t�������
�hO&���uQ� K:�0�r�$&(�@��Cp�2�oB����K��������6-�.'yX�+����̌{6��9`38�A n��9�Vl��E�Y8��۪�4q�ܓN���ɺ�3����e�
7/b�﨨��"+�U�=ņ�Y!N05��޴�U��
pg�5hAD�A�g}�J�t���qה��Aѻcq+��<%=fFdO_q��'L�FC�Rg �n��Rث��������80";t�O)A��Я�z�hr?j���E���3�©��Kl>�`kG�U��Qql���ˑV��Z3���#G��A��f����9�ѫ��c��W�j��B=�Q|1kD]���f��y�����M�JsR6u�J�8Pq'0�1�)�^�*��u=6	���V�_k����2W���̶�����(��>�Rz�gA�./�\9�z︻ ��2BJۀ�v|��PUR��y�	�ki<BOc*g#J>��}�?��m1����`�H�����<@{��X����H�~Ec"�*b����%�Q����<>�{�g��0CS�"��ې�b�j� o̲y���\�Q%�1���� �C� 5�����r�uf�.�=�'n-{�D����[~�&�7`E^������k�,0�^S��id�f���|�����W��)F}A7���+�s��7�1�!_Su��45����b����tM��U���1:�%��$�	l��7�M��W�Sy#����z�QA�AE��GK��d䉲�v!�sG�(�N��r�p�`�C�H���MdLN�p���O�ё ����'��%I�@��&P�tG&}Bˑ.ڥ�-S}���k�RĤx\�*�	x����c��x�?�vт����j'B��;?���<3�IϺyI,\q���<֡.	�:��!t r~r�5Hy4��ڧPAe�k@�K�&5dv?��_2*Pm:XI�8b0B�>�\U��C��������~�*7i�hˊD�Pn=�d$�)��ݷ�����\&��P �͐�8`d��Y!�3�`�%Cq/��_���9��\���$��B.�M~6~|P����i�������43�&L�+����ZiϬ�F��?���?`۝�hY��Z|}��#�Ȋ�{�&o�`I9R�j�y��7�WQ��@	�1��;�e�F��B��/^W��G��b���%\L��P״FB�/�;�x�~u�x�s�<I�H��n����Ǎ�}@�jm�,���]�[��.�ab���O{����T<w5�qu���U?r���|��'�d�uX웱CJ��N�Cp|�rG�����F�^T^ZvS��"a.�21� �}O�$ϼ��`��g���/�^R7��Y	�VDQ�&N�����)sqz���ޱl�����9�=�(���XHp�ҫ���;`3N	RX_?�Q*_�^f�gX0�D�r�U�%��Q������`�xSs��Y�� %Ŏ�n���jY����o_�^ԝ�]����[-�f�R�d&�p��J�y��<�؏0�(u��Ð�M��E�e�͸�Kn����`��OÔ�2�A�.��c��N��}=��!�����.����f��?T3�g0�}dQ�6�E
�[>���CV�qɔ1�8�ω%�^�D���1xg�v{�d�K�����w���0��ɑ�`9QH�̥'�;E.R@HA��:ɼȯT*�XS�e�TJ�,��Ho�r,)��4�%���$��,�wc#�<)������Ҷ�L��MI[�oa�B��u�H��L�to�6��Ǻ�O�)+���n��;����a���20�7����k��K!�Eb[���թ]�&7�k쑨�����78#��� �nA%t!���'�)��8�t����n�hJqc So�B:]�\��
�?ҙ�`I-�=IS�[ď��W�5�� �?�-K�X�����ϒ���D����i'&԰Ʈcj��J����>�Ӄ���I,�W���9ADy��G˼�I"5��|�4�r�:���f������ʳ̀��6�~V'�ǅrs�6�,$�_�m��?-�봮V�&.�@�[o�S	�d*�<�"LC�h��S�)� �wN4��{IU��0�0�@�c���/��u�,a0������/��1=�udؙؓ�*Zx@�Bh�@�G�.��J"W�I���:D��;$md���P$w�Q-�կ��x��~�������:�%_:{��m)����$<F�'73�i�}B��k
�3��?v�A�x�=_- �!�r�+1��[ jf�R�B/#�Wt�Lͼw�ԔO2^��n�PG�w�{\(��ޡ���qAh�Hl��{{���J�T5w⻺�0���)@ f�W5����qk�Tn���i��2^:�%������+��4�,��B��^N)��T׾�����t��y\汷�sYj̙��/F�v
�Bd�F��RU�l� ���ܖ�e��cT��^9jX�s�C��/+q4���X�]k�I�Z�T�Q �FV#���V���J��&�?��?�ɛ�v�y�G8iIcY_qf������o�������n11���0�k�]A��1*.���0�Y%"�>������J�P���a&PِСB������7��m';�������c��aX���$��/�]�J��� ����D�!K+�����j������ �b}[/|--���=������5�
��1��N�GR?���d/3n��J)-�*Ӻ��U:��WG���{|å��@Y�9J�(��R��;zFĮ���ЀÜ3B�k�:n�FһĆ-�W�N�Yvq!��Ϟ�]�O����v�Y�y�K���c+�kizK�B,y�_�_E��H���;�����+t�b�j+�K�WC��K`�����m/f�a~�州]Ze�S7�i�B�
%��K�O���N�=`�˫Ζ$]�����K�k��߆cA,8��;;DO�r˦�T?c��O�HdWp�e����r�����3�GW��]����Fnŏ�ݦb�T�w�0�(��T����ubh"�~]M�/ҋ�ڤ��y#^�Ae6_h�SՋ��* �F6H�H�v:���jZ��b��vX�'{���=,��_�K�6C��!ί1N~p"ԧ�W�[�<���G�D��E��I3�e�-9$gmz	G�����^e���zr�X�-L�.ј��2*�O�D���T�PX��f�]���p7>��!I��ݮ�UX4�� {��ڡ ���s����V�����E���!D��Î�|p���^�#��J�niJ��eĞ�ݔ^�hc����c\���j�@���G�:͹'�7�L����%_	2Q�dE���d�|�� U���FCa#�ٲ�vk�������oMX؝fs�O\����>� w~gE��ǣ}oe`~i�^�&��P�������G"Fy�_�:N����H�u�W�K����w�Nۼ��l�"�:H@�G�b�_�ߥ�f���Y�����t.�U���M[���G)�X��u��r�y»U�=i�V��3�;xa�|�Jx��wƂ��=e��h}�:?
/A�XM� x;�n��>0D~��|Y�������@�u-�.�g�8��4�;�����Ez���~���1�H�h�ٹ�L̿����ns�(`�e�C�Jww5��#���O�0Bk@��_��$U�ǀ���)g��N���/�
ꖅBJs}+Ò�Y��D��|T�@��� O_��4k3~�C��RU��Ov�S�Ame����y�<��QF,��T��8Zբ��5t�?�(`̀��ˎ�;fU[H���LJ�r��dOi���:;w�)%��&��.{����չq�?z0N6�@��� \y�e� ֘��t�8�'>Q�c���JWi沅u\�K�S˵^>Y�ru^��~{%夸���!� XIs�ޓ扤:1�xrB;W��x���	�qwGMP)M�7R�UU�S
ea'���oyU!
�
J��;�m@��2�G���Yѽ(�q������9C��������FƱ5>h|���0`~��T);�K�^2x4��� �8�eU��a�I�(3�l�m^,��x�B�}��c���v6f<���|r|�V�]%|���;�8"�����f �[�@<�+8 ]$9��;�qf�>Nڶ�ؒt�a��"v�W��F\.�USG	"zO��'�pN$F��Ҽ�-��I�]`&���4(h��]œ��5:=ւ
��i�@PL ����W7,��@I�*�5����_��y��#K�Ho#�*篁�E���H� 7�@�猿m�˩�k��A�F�H����.�x&�>��9�*��a�5l����~W�U��9k�\�訯
4[{���Ҩw�/� 3y #�{��|K8&,�it�y�A>H����=;z�3���>��.}�םR�c��Ҥ��G��O��h�W�$	5�[�ڵ��Cx��i��6:/��L�(fS#!4�yp�@!Qa����}Q���VOX"�<�����e���'B�8Xy���E��b����T�'���2Ix�{�e�2oWcpPX=��7�ںY�=����xK�bHY���AR�b��+rʝ��he	���{����`��;*Ta-�Z��_ߥ�	�0�N����*(�͑g�	��&8��f}�}Ѐ�3����u�HLC2�Yov�~���?��b,s��(�q����s��������ѧ=��|}��_�s�|�VP�T���"�Ju�+��1W9K{jVC��,�e��2qv��t���E�Hޙ�݆�hWt�'�p�Q	#���[y-�N�"LZ��+ه�H�k�%6��-mT)s�6��sj����*xq��'+�m4�R���CGu(L��_k��Jů�.�ľ�oFk���>o'����>��p��6q��9��(b�O[���4H\0�=��!�R7�?����'?33`���!1������%"T2s"F�t��U��&H<i^��a
�Vvv�Fe8��e�i��#m����=`Rˇ +HQS�jxW�����A3�sA1L��Q�Xg V8�-z?�' ����8ң�zCl=��q����z2�Ќ���/�� $]#Z:�f�T�o�"M�q�&�
�Ѿ��׼���EEQ�>�/a�$��e���Ib`���w.�I��#�(�=Ã���T�C���'�ܵ��E5��^a~��=(�]-A�<�_z�����<�bu�j,����I9��|n��v��KӬ�5[j���Y�}��"��܈;?���j��u�#��l7�\cΤN�䋐}�5@��ZБT�k�\���������l��f��5ȸ����|�ޖ�AgɉP��ZJk�����ZH@��*�"*�G+!L�oY�iV2��R;��W{8^�&{pBY�̟�)��c)�mQþ�b`\�&fWQ|̮r��.7o�4!�~�M�3�����A4j�w���`��<i$��m���u-M�L^�;?^��>��u~�^��������3�
i���$�����������z�3�����~��W�kNYc�ǲBg2S�d/��F���x��<�Qi�=@_�ޟ��a��rƚ�ӗ���pԉ�3a��L�Zq�F9����DO�ʋ�/kG@}jE�G?�C��i61M�"a/��Sq����ǻ��|��j}��ȳ�'B�P~�C�r�}p��{gi�6p 	�@�]c�^��)sV��I*ww.���9�OBݷ-���E\$�B��c��\a�z��M���z��"�O�8p55w�㤱�:�4P���y��!T���-
�U�ە��U] �FT4h+A�{U�
\����r�Qú1n���*^<l�W4)�@D�nEF�D�J�d�M�V��,i
�ˇI���`����j2o���Ԑ������%�@�0��Ff����U�������VF��c�n�"��ҒA9~�W��C|��a`��)%���s��]h�$o�
�P�m:�DN�~/{�ZC�|�}z���kb��\�^_���Rb��>Z����2 _�)��<��^�
�Vi#�^L��ޅe?W����ʱ�J���� �TM�s�҄ϻ��� �xpuP�T���-f4.��-��a}6M�j���r�~In��d�H^o�~E�"0ٳ�zo��1>z���g��kc��Bp�e��C�����aA��x��Y��<���
j�Z��AI*Tm���k���e��f���÷���Ma,3Z��|L���\���Ga2��qG:=�����{��"�̿	Er���\�eQ<���$zI��H�_�]�K�¼'VS|}9���ݘ��5NA����&�z��s�u6�n��+/aYJp�t�ķ� �������9j��%���h`�eGۙ���\�jHF�,�v�Q2�?����w�� X����ڄ�bR=:|us�8r��5�$��n�H�H�ਯb�#yBi�b����"$T�?���qH��Tr�L�����p����ֹ;����oh�Zz|��)�77+4C�։���ՃB�(G����1�QV����������(��'�|	�:��B�I�FP�;�^�ϕ�ݣ,�=%���X�v���nT���`��I\}[��� ì>��`��m�y+/O�e�,� X��4����~F�^߮�KA�5�p��u��'��a4����0�m��+��O�N+|���;�^_�{�
]�~���(M�M��P]x2���t1�u�"k�u���A���@mH�",7mC�}ߏ��Z-~$��K�v�(�#��7��%5��RyC�U�)������	�n�ħ��	�a�^�U[:(I5�s���ߪOW�"�`K����h�����Ӂ��g_�Zy.�7c?��Ź�#��k�@�O{ �����0���9,�IM�1ZXG�#�Iއ]��&~��ՙgTl�b,:ͮ��x���/�)\[5��A]?�ώ��fD���	gwe���ukY�L*U�3��tX�E
U�
��ﭹ zyn�{b�Bg�`���1E!r�[x;��$���g?KaOMh�6@W��mr푩;sda�jr���9j���2d�院�ŢO#j�;���!C�sӄ�N� Z�/��rRM-}T�� 2�@���@�ԴI8���5wc�7�ꘞ�WM/"��4�kg��5g�j�ݫ� e^L&�p�-�Kf�.CZ;1Z�݉�eW��(/��M�MO[႐k�t�ݒ��.\9�~rC������L�`֮����B�f1�ȁ���%�8e(Ƃ��:�	��j��@v)0S%%ҿ���� ���#�87���K�v��(��d_
�s�]Ɲ�ٚ/-��f*qh$�(:u<9�ǲ5<�_u�-)��c�RŽ66?�ϋ��6?:ܷ{6n�,nȥR���h�qSK�9o�(�R^�iqo�*{OaS=�|�GX<Z�C�_$�g�es}Hx^Σ��j;r�hX�P�6QH3G&�[��vjP��f"�y��뙂[����	7�w(�z���y�Y�06�2�Ysc]�e�G"*W�F���LwD����Dm�׳�u�t�!?������m0ڐP�Hˍ���4�d�d���Dg$�n�*Ǌ �T�Q� p%��`I[HC�8t\Y&�,���������pV��o��zH����'xj�E!D�����w�E��1�:a) ����X�����3<�6���_K+��,J�T������%�W󡷅�@����l��" ��lh6 �cȏ�<���h����Il�ϭszg��`O�&��'l�yꞱ>,%_geYؓr�T7&�i�*�L�j 목�1�M��!Q�ׅ�������y����.4_�r���G�[W�f�#�� '�wt6#���Ŷ=@�5X區:";���M��@j�߅�^&����M�M�FW�09��<�ie(Z�**����\��'��_��[K��N����j;�w��qD��*G�
!"gӣ���U㎨��;V���I{�M�������
�HeF�0	���w���W�0⒝t6�"Y�)Mإo����.o�/vƽE��/ϫaJ�
[�v������xN�L[��{��z�S�����c��/%�E�1��y}(_^����Uȉ�<m�F���J�M���WZ�Â㯅:<ʒ���@��A��ɷ��o2���nD�!m߈Ɇ��x���s�s����l�[�:�]��A�
N�� Y�R�g������D
|�+HkZ�R��$�(��AE�^��u����ހ+@_�8}d�(�r���SFӼW��e�y*��8e H�.l-��q��2�u7��(�g�!S2��EGVȤ�XNɿO&I��x����=KV��r�n�f�z�O>yä��8*lJ���x<�s��"Uqr�Ph9x낋BcWd� O��p!�8���������<1�qa��87�ph:J���	ݣ�K}�"Pf� N��F+�{�;���� wq�f��rvg+M���A��2�_���)��(t���}9Q��-��C�O�R�ݯ*�O�j�"�l���K�}�!����d�M0
��`�D�V$�>ӽ���N�&{s�SN�-���)��u���?BpX�۵�<L�[n5�H���8S�i�Z�F�� K1!��!���	���K��$��D_�:K�c�?/�Ψ۾�P%�+�:n�Lj
x�����N�6���=;�*��<�#o�,���qGG�"`��@��ki@�mY<���f�3Y�)T.}8C͊�B.�Z7cC
m�A;���F	۹��vY��!Ȕ��y�c`;�����OL���ss���"\��D��t̹/\�DR�~�,��@���%σ�l�#aU-enFZ�JأH˛Wᤦ�l�'����o��_���G����H��g�r�"�߆�i�2�>���O�X�4�̺`�l�qA4��]L+~�]���urC�-OT��cBa�"�RX�����b�6��w@���P^)�Vl�t�1X-KG���y�YF���1����@�O%05�7{��0m<6P�̯-�q%ul�є��1۱g��Zb�SqB����e=�NȨ">�a<h�.7�-u4�ʽ�+�K�7��zP�FT�8%�Iʺ���p8k����"y�p�D[źwQ0
0V=�{��ַx��sG�K���r"_�ܦ�yQ����6�֠�p�i�@+:R���S���zn���\M�ȃ�0t3ŗd�B�6�9�NB'���ٖ�_B=k����P^��┐l�y\�F�J�9D��I{�)ZP�L��ݴ��Y�P�X	��b�Q{G�d=��J�>~�x`��g�=�ks��%]��^̌rI�ܻU��v�v6�������X��Qh��F�X`���<����U%�W�c+�_\���C~2A���p�k�E,�s�̆K,�Wb����P?i;�/E����i`IzKyҸ ����
c�l����+0����q�$=Z��|v�&rc��wm^n[�wv��X��p/��{�?ѳ@.fw��Dx��c�㎍Tמ���,Y�2�ʦ�BdU^&���Pa�d�̌��U�E�\����*Eoo�)� ��Wƀ]��Q��h!V���^2��=� ��gy}�˴5k�&�
���D�
Bu�0
Q�p%i?��݊���a0❓�?DI_�Sg���
4�l4O;P6�}э>�{��8�>{ϫVrm�:�ށ<�Ṅ�|��J�̐�3��������yТsҲ�߆,{�a�Dh�?U#y��B}��]j�'Jk~��fM$Α�j�nf�}S��1x�&��������������c�4{ǥ�<�qnM/��)���1��	�9`�iAcǎܕƷ0
p,�D�O��� ā$﨡��������q���HƟ.��/-�W  XQ��-rt�)��5t>9Ktk%7*D�����TL��l3�l�֖�u�otj�@Ή�\/6RC�mhg�[��P���)��h,T 츉i�_,��LYPk���3ʚq���5�.'h�����ꡪ�s⚣�T*ri�ד�9'۶s�ȿ� F`!��:f4��Fp����Q�a���d�W,�))�����Ŷ���k��i�l0u����|n����wi�`{�a�}Jci#�2-=��*�,�kC�h*4�S�πN�#�cf�1"�Έ�����\/���vh��oG�����A�¹@�.]۔n|��?4(V���
;�=t��|���������j6��8Ty�ңH�vqQ2/n�����r��s,�/bJ�ة���V��\B��B�v6)UP��p���w����f,e
��^5�`��١񕕙�$p�Į��H���'خ#�g 6�	�M���PiO(dc��9�4��g�	3��l�P�D/����VKd2� ��n�R��0�����j=A�I�B
V���s16&�m���|�a'��S�P��w��U��o�%|�<���m��h��|��M���:,�m� 0�Q���u�Ke���n5壩ȕ��qE8����l��-���G� �n�w�k(���4Y霱���WF4�bZ��IJ�?�b\0����%G/�$�`ݪ���BK�`\��4���[��='%'7]����n^ca�H��Wۗ��8���G���]ѵBX����(f[ �D���Uo���9��Wd���X���$}��G����W��5�7�|f��w2G�P�h�`$@ڸ��S�K���yo؏��lN���]��&qS�՘�E�.0{ԙR�ս��3B��)��u�^0��0��"#�(]s��dT);��ʢr��[]���L��0ݢ�ki_�[g�o�V!�Y��3q�}���$k�3�#�ȥˆL�B���dh���B�BQ����]�p 3��B����u u�%z�e�Z%�u�_/�M����P|���o$����װڏi'�As7d���^��B�=��K�k�.�lh�bI��#���w�K|���~�u�8�$�38.�I��S�EX����@��Mw�?�J��>�n̈���-n��D~GLG�I�z�G�/=-�\�����	(����ل��yT3Mj�*�D��t���B��Ti;��=]�,C+�>Uu���I{iu�'��.["�!��%�ylR���{�3s�׬{�������&k�s��>+몲�������,�J��Y}N�cR�¦3)��m_*)��'S�!21���H���X�,Ғ��L(މ!ZQ�E�;jǸ�h���u����B�d�KM��OX���H:��τC����3R>�o�_��op��X������8������mya��{k���;X��'�n�eT������XZ�a;;��Yך��DT#�%V��f����U7�<�$Z[��U;r�L���ҢE���0�gv�:J���.��,����֋�
D�����x(����)����_M$�+�E������=M�z �6k��%��q���uX"ڏ��u��V��'���}��Z����O�Y2r2�)�0�l�E^[�r����Mlk9�������/e:�{1�k2)m����q~E�F����x�\Dvq��k:^�A�(�z������,d�r�Y�'�R9��j�e������HK���~ޡx9f�$���������݉�dA8Ξ6�AQ}�<y�i&gR̫��RMd	nz���YA��:�y��DZ5�"R�j�����u��Ӓ��,�x�m�FB�U��~DG��m`@K���V�krf����A'�d�k��H��\i��E��� ܑ(��*.?����r!�NU�e�ïe��r�EY�Dy��g-Y�����K�ua]�~~����-��҃�\ !�d�oI�^��IA5���h�`�v҅w�֖q�2�t��H�@g�u-��V#�[���,�<��u�P�ݫ����yi3���W���u#ڞø���nu�G�h��ڪ:FUʰ޼wUa()žĤ����{�T�E�dm���i8h��13e�t�ә��,�g9��1Li���Т�+��k_���+���X�i�m�n!�(�b����RH%�]޵���'�Ǚ� ]�F���#_��,Q�ͳ�u�������63�I죸i�_�3'�W �����5��?�ҳ\�S�OZ�)6.8��ЈY�'�7;��4�I���/�dE��0&辧�଴_0��v�bAٯn^S�7l����0q�t�R-�ϡԿy�2�ՐkŒb9`*
�8<}P�U��&�usN�9#I���yq<�#YR[��>���f��J~f�oLD�����Qw��KA�܌������g��W���Hɞ��븴ES�5��R��t��ƾ����
KI�TkY��O9��d��~�eՔ5r+�h?�{��s��#� �����\�4����|(�2������V�$��p�����%�� V��d�|i��F�?緬I�9:D`1w5�G�l�j��z��jsJ�L����Qwai���G��B�@7��������pZS/��Av.N"�^��E�4Q}G���b	QPiD��%���[q����{�Xs���Yq~m�!�����K�y�Z�Ac̽1�&i�E�o��`��z�JF��@{>�)%�	��TT��9|���J�����$�SVXD�VW��gF�a�͞�����oV&�� @���)s���R�h��5�("���A�ǤB�.�v��t�g�(x���Ѓ|�ɺ9�܁�Ճ@NpF0�y�;Ŕ����/�#'�chm!;���U'Zh��}
�ʀ:���? ��?Lp`1�;K�w'S�:eq�[�Jl�4R�h;W�A��d�m�L��i��?��^�݋��Ϝc�꟯v +@���C��<�E~7��k3#�>~i���8��m�P�q�e��-K�8�*����{�9q�{eO��D��@	�Q\{�r��@�EnG#q���E1����XI3��Hh�ui��3�Ͷg�wk�:P�-x}S8ќO�>�w6�-�����w�ۨ~KO�D� �XR�L���2�ӵ�U�����s�j�n1&�@��6����q��b>��<��+��#�Vn�}�@O/;�/�B��(����tov��B�YMɗ��Xg������;yʑ8�[4��?sV��Sν1H�Q��v�6ښ��|M<u��n>�,���;4�";u	�W|��Ra�-�����7����9���?W�fz������yLENc����*�����7� =d�x��i6(*1$�^3kB�#D�>���Cpn���O�!��d�f#e���Q��@�d[l�q���ɽY�J�8�n)@��&	Tx���$�I��,*�*J�MI)�`X���f�TgH2v�ɑU���l-8���b��H�8���`l�ܾ�=�ʅ���߁�s�^���3a�["P��6j:k�/�r�	��F�c�\������6Ή~ f�/�H�R�!J6*ơ�e�Y�p��FbNO���r��u��U��X1���,'|�,)��>
A��#w�V&� �旫�&�r4۷���?IAE�݁!�Z���8�<a�^�Kp�E�'3�;��;nU��DB96T��V��^��E�(�n��b1���ubv���a�i_5�I�#J)��門N��J�{�{��M �-��(��T�D��I����Q��~����6
���&�Me�v�mS��	�Y��%�e�ոWl��&z��������R�nс�!t4h$��l�;/	F"�&`~���¾o����>�^�"q�_�ƶt{! b�r%�����V���ޘ�`�J<���'�<���k9����)7�mE�
�^�Y�R��!�����X�݃O/��R(o���k��\��L�z��BqX�+$�z�Af4��d�Y|��-�C
�bɻG���P5��5�����@H!�z�̂o��1�?�����c��3�ރWv��vM�0� �(L�5���B�fņ��'�-sWb�an1|�Q>�t-Q�t{#䍂��.��� x �^}����9��u4$�
X�(O� ����m�����;(��7�y)'�V����*�f��W�dG"	a3�o]?A�r�x�4|���6V�JK�^��g��6���l�(�+D(��%:=�eO[��S5s���~JX�u'�^�>���h���"��i�d*�姦?3g��J�~5?��&��ox�����X�U����* PaxΜ�TE���(���^�c*�5g6Y��ix�Md!!7,$�3b����4�0
',�����LpTu�L��9�(��Y��
P����̅��ZI�[M۴�ʨ;/�JTE���kUȞ,d4�Ki�u�O��l?���끟��L��'���� �����s�����n����{�s���S@{Ƨ�݈�/iC$��m���a�i{,.�z>��%2�.H�����0l� �l�|��Y�hG/樆�]� ��.W���i[�+uo ЋVQ��O�ؑ.צ�`ީ|�QU��S�}F�*?S�6&�$H�z�����Vf� �P�c��K	�Q[o�����F�,I��āӈ�z��	O��l���Sp6k�JHV��Y�M�I��@�0*u>��>R����+Hg�=g�
eR�x�|4ڬL@���?9�W-��+�ѦiWOed����V3�:�),v�����v��R�wat�gޠ㫨o�@��(^#Z-'��ڵ��Q���%L��=5|�%���v�`zEZ�tM�&���%�]ty^0�����ǫ����^"y��T�l۷>��K<Ƙ ;�܌�ԍJO|F9�¹.� dk���)�`}�Q�<c�O�W��G�9�kV��7.g�"G7-�o	�Ds��K
A�-	d������:�`琤.l��K<���ԍ�!3�jz��PE��h���'$�P�IMYyBS�M�E�&�^�L��-B[�j�w��WΚ�AXb���H#��O<�t��Kpd��S�2A2�'P�o?0b�����(��bl��G|�>`�ꜥ��|عYQXJ{2(���֓�Xhw�=�B{�ݻ�D�����J]�ᙫ��>a�r͌^�� ���64^�|�����2̴R����1��G�>���l��=T�K�%@qn��G��ô�\>_o_��۽]�a�`-��_�@9~���a��o��X�aN�f����/Z����V���X���v'�\�ʑ��.��Y-� ��5�B��>5�cZ|P	�E.�B��)���l�v��a�_��Й�B��L����N ���=�>����i��MS5���S������8�����q��]yLQ�����5��ӗ`�MJ��7��YC�o��܃��F�Εni4�����\���z2�>�D����̄ ��	��S�:l
��4]Y��܅�ꬸ��C~Q7���z�g��C�t��;���v�D�{8bh��x��H��ۄ9��S��޳���
���[��Hߢ<\�}��!��6V�I�Ck�����ķ��@������u������lF�����K�����Q�4�Y2̻>P|~XO� ;�{��u�C��eR9�ó��ެ�m��5]��w9� ��	����<)�.nQ��<ģ�5O�iYzLʄ�~D�TX�g�1a���U��Ȍ�S�kgZ�.�#��XL��
�++w�����d��ձ�c.�:?Ni/�M���0�5�A  �r|
.n�*g�G��[).m�[_&Q�obUƳB�L�h���TK<[5[�)v���5�^x{�&r�
�A�R�7�O��R�i��`�2��@\<'],������y��=͝�T#4��t :�4��aR<Xr]]1��?H�T���g jM+����ح����Đ_�n�>澒��c6������4]�ҩ5�	��Hyj�sr��ߺ�-ەLg>k����n��.@t��:����Jm˰9�rV̮W�2>��b�R���:�5������y@FTS�o G�iv(f�R��`/[٢8;^뼛,���da��s���#�l��$���Q����s5,M�3E���j��� ӧq" }]n�x�Kv�#*�C�Ȥ����{�q���3�ñ�6)绨�� �2J��$��U�!���}z�i��o�
��2��D����@'�UQ΁��Q�	l����&��[���״���\���<�ʻ��x/��x*�mO�œ�c���$pU-������������`@̀�@(�׋'�������|6��z$0"�u���S�(a�ڝ�b���&r!��-��r�Ϭ�C���ʟ���C{���P�d�:�����i���/��I����HS�h<w�g0�t�P!e;�(�?����1?0y^�J�xa��c��?�>�3�[&]��ΰ	����g�,�f�Ԋ8�Z��Ag��b�j��2L*`����x<��E!�W��E@]�����8�uP������HTJ�P@)���*�4!X\-�8i5C�:"�ts�n�њ?�-�@v$����OԀ0�-|�F�I�9Wk�����s�3�̣����B��i�v�F���_77���|w����
��ǆq��O�F̝LQl�p��ʇ��^�(��#
����k�*�GX���9�5k�.�|�U�K�ܛQ[�z�R�X��FLg`��壶���W�_P7IgC?H�a�u��¡/�:#Ӷ�2���A��7{��1���	�KLW�pĊ$��_��Qu=�@�}��>
�#�NM:7*�;4J�X�y������McSl���Pv�  v�F�g����}�2Y?sc �7�i�\25�f��Z�҈Oٜw֕�qW��[����i��~ٷ7��MT��C�V3��>t�v�*϶�z���H7;�N�DyYѣ�I:�a��5�p1&�Ua���kC':;�I(֝^�#�x�H|���ۂ��OE��Ŕ��E(����OX��}3v�G��<=�D���Gw��z�d誱����g�8�Xi� _W��S<��I�?N��5#�y'!�����a��o����2;�S>�~H��gĜ1C���<W����[шre�N����#j>qWi�*�!��T	�̾�lJ�ħ�m¥5^����%�����؆2-!gd�C[e�\ ����j�[/{����^�7z..���
#D{�v�n��-@����?Zp&� ��s?�l�3��m�W��9��.���@Ɗh8G%�<pn�[��e��0C�>���|���Zƛj�O�8��R� F'm`�	������d�_��D��k���=~i��e֙,Z��FL��2�jDn3�M�Oi��&���:gc��ԕ�yj?t\�Bh��:}�'@�o/-.�4;bU�����Gӿ�(m*&��r/� g��C3DB�ެ����K���c�I��X'���ҍ˟x��{�%��T�6L� ����N�C�U�y���,i��<1^��[��y���/ K�h���k�wp���0ҪEՒ�/���\���Q#�'^��T���/KIV��p��4�]�% ��%�k�?
�#����GrX{%J��_��6�@^|�/,��%�����TI�7("�o-�*�n�K����t)�l���
��*����s<�ЂO�ex�����*7����'�X(�1�����k4��'�~�%�����*�88�5蕓Op;��A��a�����#C��k��[��o{��#�|b]f�*d8�r��>޾�I��  ��Np��ft)��}1U���'��2���ć勴_^O��Ye��L��|�Ƚ9�T�����O^V��~,.N*�#�y;�2'K޴��۴�gt-y[Ŀ2l ��G~�G��2��l�Qe 
���ma�Nc�����������S��yVl�I���7��}_O�F8��IwW
��l���@�R�uh$c+ndI��	(J���hY��U�]?�6}��A��f�\���k��~�ց0U��HO��X>)l �Te��~����ܙ.�/l�`��{�iK]�:&�1I?vt\�Rkj�C�������fE�NS4j�OM(v�A7�Iͯ1��h�l޸��9��kq�/�#����d9�}�#b�q�@2@����
���Aפͼ�QT����k��\�Lh�_"�/1@��VN��Q�K�9��l����\�3���8է>�w���~+�ڳ����QVk�k��Ei��21$a�]���q�;a_w�����+�ˎǞ�d�j�������%�i����m�j�+�kI�����%g�GF��,D���v>	�s�����P����\��*>)ǩ)�����$���K3ufY���ݩ%�ڎ-�����kF�ʄIbO���\��`�8Ӻ�����'Ճ!X�7P�8��K�{��jU�zq�C�"0̎�ʙ /��A�0#�u��$&�a8���w,�oS���7XJEW�r(�h#%!<�$���4��$�	���V��O/�]�Ch�\�S5	B���������"�;�F���'�gy{�B��AD|U�	�����aɝ���Z��(�@��
���exDg�tM�J�-�!4��̵�C;�l#l��*� j���`ρzJ|�w¸�ѭ1LC��Z�4�M�g��\��w�!�)̗����q��,ΛUG.f�$���3l?(���J�w��|��wYu|�b�����B=O���Xq	
&�ݛ��p�ո�	钮{�M�|E7��YW~�a(%����iԁ#w�F��b�X`v���D�K�������?dxq78{&{���hG�˵��#�P��.˔��zm%������2�H���V��[���[԰m�唸rJ���2��<�2O���.��j��jw-�4�P�б#왲/��XiN�)�;Gg�����|� �{o��m5��n@TAL�x��P�Q�15�����w_zX�k�����`�@��Dޥ.�%�{,tf�ќ�2ճX�V�d[��3j�x'���ZVw��8�̚H/C�Ϥ��˿�r:�HF@(�yEf��o��g��:������+0ess�zMt�w��Q���;�^Ay��-lXS��nK_$�+������C��Ѫ�i\f�0uO_<_n�U���y�����8~mQ�m&�u�Y�`Gn�<6R�{��]�5�ٍ��]D<m�j�s��nI��*aV*���"��_T�x�UH�E����Uz}��UM�>�I��h+�|)c-=.� 3�r*�=>u*�-�P�1g�,Fab�|�Ba�B�7tj��L���ͮ.�8�o��Ib�J��6�������G���ekZ�����s7�-�C��5O�f���lj�����mh�1�>���}e���=6�H���MȪ�3�������rfMX��ǂj>d�ie���	�����e�ӥbTM�
C��������ċ5t�A�`/,hZٗ�v��!p�!�4�[�1���݉��k4�<u�LL�g�M�"�\��)B�Em�g�o�綯 �TVt,8�OZ4�a(�`�������l+X�X!|(�u�vdg+�d*#,���kA�#��9jE���p}�Ѷ�MOꢫn�p��Քr��$�sG�R�:O��,��dT��M�}!]Fz�U�	'��X��8�zM�4�]��ɍ��V�J/��;縇���_Џ�V,�&�bw�#0�
��fR�����sho.p�ZMH�z[JI{@�!���(�2h�(�ٌ���o��K�����.0R��3�KO�b̪�jc�ߜ�5�g�����6F��W�5n�S�$�M��9���Wy���o���}Q���&��b��� ����D�_ǽ��
�����[V��v	13尠-�d�T��]�ϿBa0�+�����`<�+^�ZzaϚ�@�\���ܟ'�Y7�l	j��~�dӴ��، �A�]v�.Hf �P����F�J��}/#O����;�g�N�	hH�Õp_�8��ʿ�/�Lw�5%[��ع4FmC�mg��y��$uj����&\��v�G�]F�[@S�Y7�;���BC^�Sq�և(����
d�4��X���wo�^���{/�h�������_�{�~q�<�+�H����?�M1���w���y�|��h��@��}߀]��q����-q��u+��F��zxr%'<� :uǈ����h��J����k�#-�2|Gp�V�󎗇 s��ӂ�8�r�F��5؃p._�
��ĳ�@
H9�AP�I�H��/�?���7�x^lkՍh��S���=وB���������"����T���lc%n��^���c�K��@�d�b�J�d ����<S��6R�ŗ�\�E���@�9��)�.Fu|f�I���<8����Gk�z>�㺱�2�#�k��	_��|x�C��hX,�jiìV��:������brs[��������C ��.l�s�8sM��k~<ф��yFX{͟ʏ5t�r���d�[k�`bJE=?Fs(ڢ��n#�r�&�"EH�@�=�0�vv�_*���T<�����"���^�7ؑ,��N2Ko�_8�����zF�W	Y�OU!U;*H���+
m�,y*���.����[�~���Gzb�T�N�N�&��οח8�\ԑFp�z�@Gr�_�ʎ�^�M�+�&h���٬q�]\?�����N�[�˅�������K��}$ l�~c������f*��y����h����Vg�,�f/i�V�xz����6���juIj��E~&��?����%�DG�'@���R�ү����tl�	�/9����c���q��
�\�Pe������W8��2$�X������)�#�G���Q];�n��Q\F1qx�3aB�������ܾ�;���+��,M������ǿ �5������V����3�I��]�!��]�:��i[8���t�x/c!5��"ԯ9�;�'��'w����h�� D�x�1 f6P���6�
�ؾ����_J,�6c2Nl\��|�Ҍ�j$fr,j�������-k*#��ܬ�R��V�uru���{�������sv����L���U�T������=f &S���1�������b��Q��)��- �S.Yn$�
y*c��'1�҄�r�◐�j���	�̏���=Vv\�>~H����S�
���:9�I��e9liA@����Vi���h�ı�U,Es���6��A[�c�p^�^4��'���N��F��bd��/7�]^bC�0��ێ�e�^�o�ᯩ�G?;J��j�@ �y}׉(`N���p�)}������bH&c��f��f�VW�
^���vf� (��DC��Y�S�&��:G�F
-o ��I�a��yL�,�g��G���S#DL��ǔ��N&Ii������X��V����=IV���o�e1�P��Y�L��i_��4�o� ���S�__`�sup3�C��Ơ�F�����%����l�͎�ͥ�fbn|_���N�S���i!��x���ц��Y_���G�~B����9Ů+[�@�x<��u�T7�ĝ��'��-D>�V8|ޫi��3�p��$����R<V����,)��C�E�$̲1��L���*,��27�(8�r��x���`օv�R$(����I�o�8?}&q� �ܾ��
��٘�; =��iU^����ΌZ��^���* �y@E�m�g`�L�����3+e�7,�Y��Ġ�/
-6.��X��Ո��7����h!8l�s����"�}�z`�ʸ�f��^ٓ����K�� <7O)�lw5`JR�ͨ��z'x�<<����
@N�S^��b��w[-%5F�`�S_�a�^-�D<�_�T�"o� ��$�7��y�_��em@o�����(?_� �C����2�x�R4p�]�E�:+=T��#�3�*v(C��H!R���i�ԙ�yO���K�~*��HdR���~� �Ҽ��S�V�a�>��-_��-W:�������y��)���n�'��]*Z�t���;�[��q@i�d�Ԥ� ��Z�z�;D��U2���j.%Y��V7�c��6_���!�/�[�#bQ7� �b�c~�e�Y����65
�=o���v#�ca����&�m���1�R?�z~��NH]�pY+��qKO:\Q�!�ddC��`�*��6�p�dL�X��X�7ץ��ud��_�=@w��Ai}\ ��{k�A'U��~k����:1y���F������\0ӧ��a�vO˻'���Р��0�� ��dw$j�v� R�k�t��F�Rl��D�U$.=M"i��P���2(�߅���V-�������]�l�x�����i��Ӭ��o��6�I'q��������|h+b!7�AA>GN�|H�da���os��J���(��`�9�	��=��h@Y��oHRh�]dj���k�Xl��܀"�����i8˵�;2�!�#C[Q��ا�w"<�ӭ���l1�!�A�����r��#1�����o�⤛�g�o�%/Z�O<~�~^;.�����W����O��<z��|.��R`iK��=0����y��ʀ��5�ڕ���iPD�F<��Uޮ�l��?�Bn2W�F�9x��v{�G|��*8�oC��n���+:�n�]�2g�#s�$��Ɛ��5�kIy}[ǈ�'J��`c �x��+w+W����1X��vtf6����e�5���'��O��xK�,��]ŨE��J��6
+y4��cS\��_F���^n�@~IH��~��45<b�¿���*	[�IA�~�f24"DB�́�}@~1� {�WMB�+\�1�Q%�kÝ�ۄ�����5}b�K���]G7J#�*��u�(8$,޺�"}��h��_6w3r%����8M��տ-�q���P��+++tn�KB�o�キ.ג�B�n3�y~Hr�.]�@�J1��&U)40z����}��L���B�Ϙ�?n�x�]�&U`�{.�I1�(�}gX��I�ua/R���>rNGyx����l3\N$�j���.8Wq��z۬���gK-�4�>%�V�>���rg�u�(b�K +��s��0\��GG���o(_���.�%�oށR�]JK:j����wQ��1ƅ}�c/�~-��(O�y�MW+"N g-+"��B��ɨn�b-�#2� �:��6�T�k.|��Լ���3i����V1;�|^����Ͷ�7w	ù���K�u����7��z�{Й Aj�[����F6���i:&��s�#U�f�֣K/ƻ��~(���Aݐ���d����{����l3��5�Km�X�ǌ$$��䏨��)��Y�E�
G%��X2��$���&i�)��}�k�N��q�W�*+Đ~�r���]��D�@
ٛ�CĒ��j>��c� �ȉy�РycOd�-����%է}6-� �bݡ�g��� �H��%�Z8Y�[�[��o+P���9���TO9H��s3�T�+B�g�g��	s6p��@e�S�k59!��ǲ�?�)���R�j4�9�i3�o#P/N��8
m9��Տ�zX�!�w�7_�g!찆����5���Ҵ�l%6W�=�xY�l��/-e^�"^>��z��^���$��z��P�	�%s� ��x��j���]G"���¹�6�#8�T�*��0�!�4��[�1ϯ���������$8�|�J� m�_��asVt���-,�b���ax��$V(�����-؉L�l�L���c���q$��X�K���=����8���5�
ծX��v��Xp"?���a=֢��h��f@���y�O� �
0���o�%?����	^�+�߻Q��Ҟ��ٚ(�r0{�d"i��[Խ+M��_+A�<�� ݕ�yNrwɻ԰����$Z�P��a�7��A'���p����ET��s���:�i%9���[�9��:�v�����	��z�i
m�۩�E[�\���	螲����.��ۂx;UbH���,��i�o`��v_QWhH��`x�G��A�4�n9�j�녹�M�^��dᷤF#Ԍ��I�`{��a&.�g�Bo�d��@Z�P�cZj��_�m3�"~���g�f��c�p8o��c�#q^�D�zM���f)Bd�~���ʻ6S~n�0��iНz}�!*h�ٜ}�f3a�7����G�����Ӽ��̥�A��<�N��J��%�u��~����w�!s:\RT<� �3���Q�hw�A�")x ��%m��J�q���ո_�R)]����U+C��\2�@P)A�k���Tڃdc�g�DK�����L��>�q<���������^S�޵�����5%I�G8��olP���]]y$	:?���1Q͇�2�EҢپ���ε%��=�\��aϞ@���4lP��b����a���گj=ן`w��i�@SZ[vR�Ey �a�9z�Jp�nZ� ]����`YD��5_�c�T;Q�vxP����p��	 +�KsE �F:��YE}��k|�s.d��	Dլ�o����������f���@�vXR��o���F$u���C7'�:U�vI�[��r����/�2],$$��ke���c����Ӎ�AV�Y��n�0+��Ē�N�O����xG�[����G�O-��Zo��z�i�	�)���G�I��?s!�N8�����y6��v�Yy�|�����I����4W�9"1�/���Cق�	�G�DpR�>������)F�U�9�
ې��jhV��]����~��).#�*Ca����s��E�_�#1�7�>ix�N��{��Y��x0���1����K�b���+�I��{�b�G�gp̠�e��&>��n�>99ܹ4����'�9t�j[��wv\� F���]Q?�tU�N�T��}�Y
��HՒ��C�bO����t*5ëo��.i�.{���s��B�Xr�? y�#tSg�
��y���lqU�6��YE*��?��HܘEUf�kc�5�8N����#;��G�E�⛽k:T�,�4���-v�*[m}��"���=�3��I� ��P1��?)�o4�
$1�A���y��d�@	���Ô�؛o�H����oQeǬ��BP�"%�;�3X|�粒|q���p����N��Izy��`m����/Z����҂�z<Ҕ��,�[�I��H�ſ�i -}����!�+�c[�A_Z�錸�d6�.��9T;��v�0�`YH��/Cd���9S-ؒ����f�@���`Ĉ�9���c�3���W���=G�3��x�5�EV���.�Q��&�K�n������#�s���!�_�%�F܆g>��#aқcTJ1qPai~����N��+��gݡH�|�(�[�|ןl���k������ ���ecu���`\8!����>���A���;H���3z��JMMk7��O�eƮ��_�	x[���i��l�eT�:�7�Z�$�*!��;E9�d�q��b���	��zL��'}�8���Ȇ�ǡ<�$������C��rg�y�+��l��:X��>�����  u���D�CGĺ�7h(l6���_V���Y���MH0��:����7�[:�ɫ�{�T�>�)�ٹϘ\�$�cr���B飑=�A�E���֏�n���P�~cM��������A�{&[�j�]�t��;�t����QZD���l�6}�w�w�F�݆��T!M�p!�����f5Dm.�����5l@j%�m�o�g����g�#����z�l�x0�RG������"��h��$�k���5VdqyT����*=�}��ɠ��d����2{ǯ!o��z�n>}�p�I��w����{�*�e���j`��{Y�_W!��u��JGG�jNe�lC��@N@��t���l1�ڸ���|'��;����[����&E�2w�XH�Ihl����\9��p�j�G��۔�@Y*먏��6n��2Zl�&��~,�!��|t�M�%�'�>Ã�?R�u.�О���u�K�R����O�I��#�{�Z6�sH��;J��0A9�p�x�v���Gr�����&��i8�S�@t��%�'�]�ؘ�'q7�4e���u\aJ�zX�ûqݰ��(�/w�M���z����@O-0?m��T~f�.�|Q����OB�CGFs�d)Z�ɭ2Z�)Z�D�3M>�>q᡺N)Fׄ5s�] �2&]d���������R�H��r�)��(_���ծ.�)��iD�KYY4�%8���*��sH�	�{H@��n���)0���/<��#VJ�2r����D�u��+��N��Ԕb"����U����}���׃�(YH�L�(=���t� J�n��=�=z��/�n��n�O�G��
����v1#7�IҜC��&߸W6z'x6���+���AG��g��������7��	����3L̴]�(��;TɲO�};�U1����wp��5Ks�N�R��q㸑���}��/����NSn)U�dyw?�A��ںA�ޯ9/� �Z�,bk*����+V�/~�C��Yxp�z�i������)k�_t	�D5��nέ��"�\�����xj|��^Ԫ(8o�b��cD�fГD�������.b�Ss�H�Kjy���i��,Cm#�!��j1�/^��ƧB�B�o�����]���*�ܴ�|�{LTK����6�W-��_
@��j�ye��U/��A/h̐�� hb��ڠ��O�LJ(t�g<����]D����E�Пw�A;/�xG�G�F�4�t�g�\�1�,K �s*�%Ć��<q�Cu��B?z	�ck	=��˷kZ]���� LS�e��F{k-�&�v�&\�oc._��$��T�;M;5��W�E��5"���Y�v|��]d_��Nv����e����u�5��@~	m��
]
X��v]7b�{�Ǘ�����hh�_��E>����n�W�{)U�\N�o\5<���w} �I-0��<=�>���A͜�h&8�Z�i<�3�ʫ��������X�J�eC�8���&GB������F��h>��E���rG�NQ�Y;t<m�u]�Pʊ�K�ri+3��/�Y�n�e�����,ȑ��y���e�F�@���9����9��k�0�I6HX�Ό9�{d��˒�䂑�Ha����vZ�~��+T)�pr�&�u%�6�\3�����(���/��{��&�
5	B�O[B���⣴�3����l��WiV�zp��3c��J%�\�W�>��c�#<Da� Ũ�s�w��B�p�>"�ҽ7�<9�й��t�F���3�	s�\�x�ڰ�++��R���Ѣs�ۉ�i��2iT�M'_�z��5U|�N���iz����vN��P�C���M�5����S�'5�b#�	�[�o^���+���>��E�I���e.�(���[�"uS6�K���ȕ8�3�v�i_��8�. ̧�0l�F����j�]��N��L��Zx �V��H�E�z��=��@��yL�
Z]2��SЌ;��%��J����wZe����LA��-k�����iIo�at ��f>
>v6:�si�Y�t*�~u掰��~ne�K�s��s��������4�fNO��;B{�s���0?B� w�X-���S�XZ�6�h�6?�����j��(�n�����Y|�����+y��83�E~� �X��e�Z�>|��Nc�dY���	T��/�"���\�׆���p-�I��"S����T�n��	�e�*R'}C�|J���?#�&(5Z��M���{��/9$!VB�����LCz��2P2��z"G�3թ�l$4�T���F=�o���.�S��5�TN�R�Z���Щ�*�k̇�ݕ:d��,���GZw[����8�����&��7��kwJ�F�5x�e�9�ny��E��`����)U���TV�����6#'�sm~��:s�<��1��nl0��͋�z��f5�����Qˮ����9�xa_L�[.<o���т ]n	�r�3Q9��$�s#�%�G�H��m�{8�g\�7�mV���	b
E�!y���a�T���^z�J"�<U�~�J�Y���9��`����U�(��Z��`��9\\G7G�okҧ~ěU��E�4��c�{�Hi$6͎��_D��ũ'uY��I�T����er 
���ļ*���a��=2�~��T�e����o��of���o	����8��g�T��d�%йV/iy��d[z��^u@��|��
Q>o5(?[�*A�`��k�v�T�3���V
[R�r	=ln5m��'�/^��Z�O����6��G��5���Q9-����d�	 �ؒ��E�
JoE�l�_t5l��b�z9s=n�lT�4X���}{�9���f遲-Y��ټC�zO6��m�^��K�:�7?����?��ݶT�L�T��O1�2��!R<��j�v4E�{h�X'��&0 ���t� kn6*�r(�����E7�8u���
sӻ�;6�|/��	�:H���C�q�v�O�_�i�[�������Lb�P����S���LթY'�+NVߨ�(�(�g��z�I���=��^�'Z���}����P*�<�Y��#���> �]�$,ю�C�3+���́�2��|Z�����&�����s��}�)[�Ɏ�)P\-M�rʓϸ��3Yq�/0�j�r8X;�{Ɵ]�E�������0]��ش�B�UKqE��U��I����-較3�o���x�2.�A��n���#�0�L� -%���p�K���-�|&K%�N��F���:�HO������zi̱E���dQ0̬4Nz�0��f*E���,�
'��]�j&8�-n��sy��E���B��`Gk�{b�"�����	F���X�AӏR���b�S���ܚ��1���g����@As�<��$Ù�u?I�]k� �)����qE\��_<�<�����'�_̍�>����7��rk��k����pG~��*�/�=�J�l��pT��Z[�[�\Z��lo���o\Ő��O�(���(���b�_G�s�g��㦮#��1\]+8#%;��-�c�Ŕi&����V����V��x�]b�^0���d3����A$+>7Qȳ�`��g9E�ۉ�K)�*�[�N��BPu$�N�?m����pjz-"cW?®��/��?Lf�U�Rbq��%�'��:B�o��gj�2��%[���In���:���ܼ� s�]pF� ��#I��Kw���1F��7=��L��b��>͂�!�Ss��	�~�S�8y�ey?s-�吵�<�@R��Y��iq_�ICu�j�[_��}h'�
�PK�Џm]Wq��#�/=���l,+�ٛ��`�k6&COc\�t*#-h�H�C6k�x����3P�߇���a�n�#�4�9#�]P�DJm������B�)Q�s�9��Q�r��u?u%+s�>o�f�=.~�>�^6]����E����b�6��Q�z��a|X�&�c�2]��]0��ډi�j���5�x!�;�s��w&T�$;�&U6��X%��F"����)J�%��laI� ��WI���U��ޝ6�#şI�b�.�Da΅���������s ��:������w�Y4�M9-a�cW�O��H6�y�g0���M�h}e����>˔i���u3O_-�'�r'���ʘr�<"�RMZ20���%-W0᫁.�p�9�:D���[�wV�w�EVVpf�4H�$�jma��n���7O���V$Rf	���ыu�5l�>�Rp!�/Ѧ�Ch�h2�J���-���W7W�ܱ{
�OHŕm��[:6�@�2,��H��!]���W���CF�2kZD���;B'YX��W�He>ˉ=�s�ԋ�D�r\�=x%��rѱ'v�"��E���cZ���"s:��,�B�۫��*[����*������>"��B�xO ���y�]⭽I^HHn�ۿ���D���>�� ʨ��;
�4n���ޗ�j�,ա�e߀0r
�O������{
N�v�#s�V�_�o�P�Z��^�׵~��knRP�f9�U��j��^)�6c9��ɳu�HLzBh��J:���q4o�������������,�jZ��$pi�0 ���ߙ>)Q��@��f]S�
Y��fx�t$L:w�� �jH$��q{w��_�Ò��������v�Ejm��|pdX5��u�ܺ�sqsDN���g8N���.�����X�%g�S&V^>Ⱥ\޳~�iax ������J�˖����D�����N�`�l��>����]���=�~���l�煈/y���O�n�(?4�0v�2_�t=���n�����N�+�V+M�77���Ɋ��
Sx�.������~#Q��s�_��7h+�G����`�}`Xf���`��Yruc�!��~�+�W��睬3�x&{���y��V��[%6{D���q�z%�H��ɍ7�g��B�Vm������l�9�P�H꾶stֱd:�bD2�T���j��-F9IC>�&��(�y.כY�5q:p���gx�$6��L��~q���m��0Kd.\�R5��ҽ�"�;���X�G�����E�����k����<xB��z��z&�4�km�[|�2�=n�=(�t^�Cn�v������E��A��A*kj8V���)��˛?���E����q�U� ���#� *��NZv�f��83Ko��
����|��.�� ��2�-�Z���������|�ƌ�s�~>��|@i�hl͖q�+�h�����˭|w�M"��@���8�X;e��D��p��H�����=~������u$�P����y��T��#2,�g����gC!����B�����5V���iN�?������U�#�Ժ���UL����)x�po���udL��o�ua���6���X��H��e���$��@@�l�e���C`��J	Y�A�MOq׷(bp��'���",���k������L�-
�亣���JN=�>J��t��"O�չ�g]VK�]�{������k�"1��Um�:�d�W3V��1�����0����|��>�"��[V��n��T;�
��{5� �-�|_gcʮ���:h:v��F(¡vM���ƌQZ����K�
'�"{X`щ��'#�c^�ǇrYVW��-s�Z�����гv)�����h�(�.��Y����c|1~�S-��h�k4��%�:��e��N�e���2?�
ϼ�J�L�}���D��e��>���:��z���c�qy�H����͌��B��1��,*_���bvn�,����и�
d���t��� ���X��$�ނٓ:�O�)�T�"��Κ|j��xd�p��`�Qo��u!��{g��#..s�Khp?�r�+\��wQV��OG��x�rG�)����aq���ܸ`|�uM�����RSe~��pQOd�
��>Y�9��g,���5X�EW��5(���?�ϋ>�׷�
�#�����
=VN"ʢ��$���t�l�fOd�[�s(���R�=j��#GvD���m��dT^�t�vͫ��@~���u-�ܝ�-�.�I�����$���"��y�;}BZ�(�5�g��"�4��\xH��b�b��B��kٳ����V?IFCB����Z������ګ�1S����%�Z�H�U��	r����p�& לDђ��Vw�?wΗ�2Ft��t8�z����8��a�k7ޥ�"�K��9:7����Ɏ��H�����n���֘�{)�1���-�cq�YR��Q+�Q�p�D����iw���%I�N�P�,lq� ن��4ZKtk�Z�ް���7GSh.<�y�u��	g㇀=*{�����mұ~��+�+����}' >W+̴�������BU�����3��S����p钫���g�
��7&��ĝ�0�_�'�O���$��}rlq���;��H�:0��)S}����N���OHL]�_����ֺPс�GW�q?�h����I�^*Yq9�T�4�Y���XMI�oEW�b]���� ^�o��կf�jR�������1��,���0�]t{���R�=����Y4~%�_��,����NO`

x9�b���Zz�"��n��h����K�'��}�Q���6�?x���&�揁8� ���������Όu��f�LM�rY_�ɉ��ŵ�mP��({>����O�V�A^�6����L?nK��/�g/V4�E%�2�S��"��k�}�~�y��V[��eA�g�c��{+�>XV:�P�k/�����wk�Sr�q�S��z��G�ƙ����4�ر��L�3_}[��'xM��.)lϽ�^Y	��}0�Y%�
jod�[*?��ur�ˬe5��f֮	����Q��"��{|	�Gcf��n�7�s13UI��@^����绲���K8{wň�"�-ؕ�by�Wc's����k��A��Hl�7�� �_D��+̖���G�D�MN�'�8�f��|z�#3�qZ�O��D�Q�[�B�^�,'�����@6;[�����3i$qg��.{���ѩE"�Tpj$j]�����^��Q��&Ǣ��ʺ�����9ϑko��}�9�iכV2��,[�y����4�e�ylA���Y�VK%�s����=Z�[���|@s�~�r��Xr��&\J�>;,���e֭��eT��������K��]���㔆\�P6LR���2�xi������g�m��@�p��gC����N��0C�/�fe>#o���|���}h�`�,��{s���� ��t­�W`z�˝�:��zT'�%��WH(9��C�0ѷ�.��l���ݻ�D�d1I��}��#rv��`��ۈv���g<k�A�9���{R��"29�M��5��K��_ǟFĽ�1ӫ�8ΐ�wM5[����n����v��La��Z��NK9,����9�Ep�i���#C� @[���%u�����v��8�9ZhFI�:��`�%qc�8��DT���ɧvxȝ'S:(9Yv:'��}���� ;vk7i���#̽��C?CI�H����*��6�%�#��D-�p�� �У��{L��v#��q5�C�>���#�z���?�	����-=��b|�Fk7^�<�ݻ��TXK�LK���&�ٱu !�����@<�r9�9 ܁DI�>�Kq!710,Un�'v���&��~�.;r�B�b^���{P?�x�i+�A�G�f@ǐ4�M�|m�N�����4\�(�r���N�jG'���۷<A��b����N���z".��[�MY D��<YfW��e?��k�������zrύY�B �Q[h�x�����U�>"��@e�I�6���5�խ(�vZ�ʽ�H��H4M:D0e�dS�G-0�y��[]���l�,�_�-l 8����P�A	�h�wKE�tiP[�m�<�h����nK�ѷ���D��0��iͩ�<���D��Y-<����.�-S�\���=���k��[	�r,x��\T���V��Qg��Z�V���i�6�l�ahFU��%�6�tqH�r?��t�v|	�^YS�˪f���H���cT��Ӻl)��H)'��I09cqА�q�W������s����>��%5��`n~���;�斶z������բ\|�0Wh�P
�����g��g�_�(47W�8Wb"�:Kzl�^����?t�+�P���<5����o���40�!Hs�@��{���h;�gӚe�7*[`��~ݯ�V!8"��'�#6�C�ѵwF���Ngm��� �{y��6�C�(Gܨ�c-BI�(�"Su{�9Нޕ���ߩ����{g�B2FnH�}��T���Gh�>JP�m�C���`	���̯�4RJ��$�-<s���K�}y��iFF�_��I��[�=������By��񜈉�E�N��B�d�=
@v�&H�#�s�O��+��R�1�T�`䝻�d˓d�����a��P���Y�~`5�|K�Ӕi㰲� �uNn#��ٯE�N��>�S�c.�������h�N�b�cW�I+�$�盪 O/�(�wG�R��N�9�'�b�����U7(l����0���X���Ѳ	��-�tO[ mٖ�`]6ܗH\D>y7Q
�v^�:`��Xb�-�ee3���f#�;?[���C�p:�t}�f��o��=�F��?�-z��"q�&������y9T�W��'v|��)�H1;��u��dH(3��sS��+V>�Q���m�ES[!g�Z,S�)�M����#̃_�R��-��6ԌJ �g����]��M�Y�>V������/�.������"#��}��*a���-� �J���b`�������uY�|��*� [%p�g%���~G�.XՀ����-���l�8H ���VY" ���|.�92J������B��L�]ͤ�^���sV�D��VG}WI˅�$�틾p�u��dCg�jf�l������x�����9{})<����Ԧ��ё���(;��lB�������ZXg�;VC��E2K���Y(��t�F
�$�R9��P�dQ*�r��nwjoQJޚmS�Xr��C��c#�5���d��������e�O�CS��XH� � fӢ�����V���%.�,C���������M��h]�@�f��!7��0 �f]I��٢J�(�f��pL�!�iv��[`e�#��G��oR�i3�%��˝�2�\�;X�� h���MOٱ��6	�P'K6=*`-�����~��>d�W�iɑL�冘�2�kO2���
�x�NKG$�3�!SFQ| �{P��� BS��`vx��1�^,FL}���O�����e��كW�ߥ�9�\8�*}�u�,�i�rT|P.i������˒�_|gӽz��C͉��sP��l��C�0�\I}� �q�'�q�[ .���#*�&N41F$�s�C�8�։1H���"qc����BP�UN�Iy1*b�6�īuk0[���4
����� �9�r3��I�U�B�=�a%R4���$Ѽn�8�p���\�q���}-�x��
�ҽfwA��Gܷ�
@�'��Ol��C�y�x�_��Dk�?6�(Y��š�~�S��s.�n���UMc�ED�n�YD՚�cN�4�Kpt+0�Z��,L�(Q'I���sA�D&t�x����l4Q��Lflo�;�Bd��z�kFY:��F-P��E@�d�hf���e�x`ۿ)d��,��k&�����-�͵���R�k51J#=���X[YjZ�K˼wO�V.�	>nx�-x,r4ؗ��Xd��5��p�A0V_�E���{�z��kh;�OloA8[0����:�6�z�PY�
�[D�*W&���,@��/�t�i31����Ґ��F�D<��i��G��¦it�H)'�6 ���)�˔?��|ĺ��~H���G���~�%N�X#��-����s}��׵
�c��@h��O�GN������Xͧ���Աf�G�+^e�Y�Q��;�Y4�e�p5)b�A c���ѵ�)�A��khx_��É��Χ3 �^��^kf�s4Uw̡���0*�:7������v��$��_2�
����*}{S�����)����C����Lџ>���:�s��)ys�3��C5N"�h'8Zk�R3�e�Lu����Ko4�ُ�8�I���L�x�r��E�OS��1�gjC��!�� >��I�fP���޿��.�r����S7e���x��J����S�Tfs�t4�����1
�lW~����0����]����8d�a��Ew��8rpuw��~�U����6��j)���w%�,����Ev�F�ű��iH��!� !,�w�Ե�x<�1��-b�RO�u�\��ocϐ7�K�dq�%�c��MD7n�6[����t�*�_H�#Ѹ�n��Zۉ`	��e�\���8/���X��ǴoȀ!^�3���(�v�% 4ʿ� �&��)�	����S�N|\^n�K*�F_������ADrMT��]��f��� q��_`bZHO����bg.����}3�Bs��L�T�b�z�L�bgĜ-����m���r�
<0޳�0Q�I|g�ƣ0X6����T�IcVF$ҵ�U����җ>�����*`&>Z*��sP��=�ҲL�S�~�"zaup�0��I5��2RD�x$�� ������\-�~rPU�b4����Ｑ�?$�����^���\��v��P�Vt��5��x"yP�(��Q -¢/n�g�q�F�����zm`dI,�kO#U�W�f�%}l&n�l��"� .uM|oFZ�j�����%xJE��
�����tH��w��ٰ6�83�Pu����7e���)�Wl�uJ�2�[q9�M㌳��%�T542�l=F���[,Hɳ���V:ex�����Z?�����a�7�G�eq+�#��3mp)���Z��"h�-�� P�w�6��A���S��ڥ
]8t�it^{Ǻ���;����fP�/4�Ἶ�=W�����b�p?\�5�le�M��N����h��ûzۖ��?u�_��*����s�y#2�J���)���1֭*� Y�������J#7�����Ue���6��l����.��ּ��]k=����u)���(Y�|bde2��|����a���km\{$�=��د/�rQ]���=�6C�A����/hp9}v�g(�)T��)�]�-�j�`�"���kz �S�BФ�1
�D�ҙ�ݢ7^|.f���r�����Ѩ�QӁ�?��PS�S����������F"&�<b�����mXҍI��n���|^��$Km���S����3<����!ߪ�//�k@ٳʂ��r���6Ao'�ى9Ւ����;�(�__�A�Fz�=v�!ҩN��!0{��C��_%�	۳Z}��V�8��Ha�A�4��jf�5�\��pej��o��iwʀ��Z&���0�,5���,ȃ��-����>��ן!��Sy`*8c.��eH�6������D>�9b��L��tm�P_�[)��y+��~e�7Cݴj�-��E]��󽂼Y�}w�T�w]��
u"Y�ŲN#k�PR	��>8Q�;;��_�~^V�5�q�Sd-j��|:
kj����bWE��ژ����ƃ0�j���?u^凅��PM9�r��ű�����,9@X]?��u���a^r�XP����`�[Q��R������z�䲉����3[�P\�@@����F��EbT������aUk�S)X�7)}���6Ǿ{�PB]��̬�*�y��S���%� 9�ɚCW����c��y+�'r�RF�� ܴ,�j2%ϛ�0٥��z�>��{�Q2��f�W�I�@K�o~������2~J�q��ƱS��������J��Iܷ9r�O�������(�3��C�dh��Dh#��I�F-�8b�
�����7�$���Hd)X���mW��%|�g��o�HôjU���lm��#����k>Uܧ�8\:_� t�+!XS�2��T_|!K��.��NS#N�`�cB���iI�&����CK�Bx��B�~Zں�^BJ���R��o�7�y���o�[7�"�.���X�n!i���2�@I咫o��M��ӥ�RB��U���M�Ͳ' :}������y��#��:fvn���s6^f�"����$f��[�.�,)����R�T��-U�꾫!l�j�v�}�h(�k��-��T���q=��������V-Je����yꮥ��� �HR����f��+�����nO4ƻ!��R����/�t�Ȋ$|�3U��9���w^G�ًG�OeXw��L�M��uw*d�EP/�������,�rzy��$]���^ivi�ɞ���.�A)��©؋�5.6\O�T���G��  �x�L�/mk��{�r��2N'E����b�yE�15�d�(��4��a1qj�O3��RP���r���d&,������^z��=�����c6,��#��vz�P��:^��\V���J��ڮ8<S�~�WB	ź�L�9�Z�|���3�y��ݻi�<���	�oAq�/�6�	b�<�C���"o�4H2.��x�����`�aD4���9�b3<���?���C ��ƴ�3�	�/&x~��X�\��*��x��@���`{�a�[s��i1�o�ǖϦT�`a���-�h	-kǵ���pA܈���X!RN�u�Q���GıʱHdw$nU���$g(X�??%��ޤ��p?�x�>�4օ��q�p�+�s^St�/��=};����q@�$��}���������21{U�����do5_����ZR���J���m��9σgJBolu��5�b��k�t@h���})6���T`�BC�2W6˼�z�e�>_��~�cEy�`l��&�h��}�ʽ�s�2��(a�Ie��$){��<?���w���2��N��x�ʡ�pܴ���Zy��<���m*5�\��@!��;q��#T�$b������ڦt!7�V��9ݵ��(3{!���8���0�ix�=�Lb6�~��Ʋ��V��|�s���&{ h(��.��5OȜw�ڏ�_��j^���+@ɸ2ן��4�ݙ˞K���@ѣ~xB�Aj��+��F�h����Zҹ�@��"�p�Qd!q;#{��6��7��۲7�R(�u�ޔ+
ewTr.~�;o�OS�����Y��Ya�K\K;��ud���'ƍ�EieS+�r�3LP�,x#7W��kD_���  XD���e�+��9��(�ܳ�ӑ��Y�>W��Լ�#�cf�ř؊K�<Գٶ�v� �
�v��X�jd������R��[ԫ�5	'oP������?�#�4]����Vl�aA?��g˄t%�U��To�3�k�t&b��W����%�]l>(�m����Y�r*��Z`a�\Y���k�r��0_,�`��f��e�����]���C(�8�|�n�fG2�|�3��v�kV���|oc��l}�EH��>�����V�O<ݒZ����,���̗w�$Z1zI+F1{Xm��������N�q�W������Lk6�[G(��1��h�j��9�my�kO�]Z��!^-�G�&��ɛ,ىv��P��t��/-]3KSP��yo_����L͡4�v�)5��y�&��oJ�g��j?&���K�	G�qn��M`���R���5݆Gjb:�Y��-s�[�6u��� inŒ�i�RJtۍa���8B���s�>��W�¥j��|Nx���ߞ��;�j;�\�h/�ä�����,x�����G
[��?�a����I
�~8q{�Ő!����=@�K��n%��mRWS<���j@u*'_�{{ߓ.VB�� *D��=l���u'�D�'�S��e�')+��h9]]J;��sdu�d�݊�1[^ZjdA�M�o���g�5�����Ɉ.k 	*Y��<�?�R՘	�>����=���i^�p䲃1��9Ms�T��"�Uw���L�8��r��n �wdȗ���z����S7�����88J�̘"�EH�����_�t�u��E�d}��ܭ��%��9��?������E�z>�T���r���#�ra�`^����	����N#Ma�y��Y����!��uΫ���������LS��l"�^��9:@y�9��Pl�=��.������d�1x�a�b��� �+�g�TuK�nn-��-\�����n>�PD���5j� b����r7<�0��c�X�/T���Q��E�c �{�lo�`�/6H����U(���j����ǒ7i�}���u�/�6��	��v�G���K仚�Fq�Y�9y�>��<����)�C���î&/��� ���,M 0~�ُ�Ba�#�3�O/�iC�dk�D�\,z��ߘ���gs7�8]R�p�4��_jMtp'z'�����/Y711�4�V \�1���H���EZ� <X�
���׌Kc��{��e�ND�5�ܿ�ͪ��r���_�O�Iʁ�y���ۙ�������(�<��8���^0��v�Q+�f�+6�k g �5���m�E�M_W�$�}�M=]R�]�h��9$��Fyd���e���{�j�{n�g��a�w����m�b�ur�W~�}^������y|�^��:U���i
�����1��6�wv��h�!��e*�zJ�� ή~�4�pM����i��v�v������HI϶����K&<��CvBg����|�#����_�zL���r=J�d(��6FݼZBT�S�1L�Tg��]���� �dA��� x#56+`�.����Bې+�x;�w��l���l�ϛ7]@��M4�����gΑ�J��ϸ��f�з����)Jŋ4y�����.�6k��87�#G�歌�亜*vGWXٓ��Ɓ�j}zh�L[�ǡ����`�Ֆ���B1)|!%$'��^|R��F}H������wn1N����|h����R�Fpn�g���z<�;)���󫤔Ѓ���<�Q�˵&O��#������9U'� Y�NN�J�JF�92�N�yQ
�{�z��ͫ��x��V���U��K_�hBێ��O�$w���ul�Ov���
B'�� m�V�H�t`��kڧ���?�ӡ�]�@�*�ss��4�(Ҽu�Ӆ�o����$<���}�;sw����!�-�W9L-�Ay�t0|~12����t^�5�O��sHo��=�)���\}�֏��/s�"�VE�E���J��<f
Wԡ$a	u��	S��L�F(Ta(��Xi��d�c�O�,Y��3�o��X�/#���948A�10H���Rx�ǉ`1ZQ���H)�$*q8b���=;�Џ���/����3ʿ�l4���I8Q��KK����G�t[�PQ\8��;aV�9٩?a��iz��Ȃ���	*��ܓ�$~$ꛮ�Q}G��<K��J�p����C�t$CjVSܑ��	~��}�{�E��fH�xNx���sY[k��^�`�� ��{yj�sK�;A��V	a/��iz�$�T h�C�
؂󠖩W!�-�d|��e���0��-������O4�)@��!S�� �=zՖK���*�i�۴�Ǜ�e��?���׳e=n���w�����{�^�Ԗ��0�S����-����o	s�B"��ݏE��5u������� Շʑot��]0��h)�GOH���T�{C��C �6c��(g���y;I46�Э�}���"ɛ�i~^o9�̀���;�hlE��)����ԿK�5-�Z`�)<�C0�{��c�W=kOip�w:���Q��@4�ҡ �ZR���^�$U���9��%����u;�o�&~T�o�gU���` D�!	���$"����]�օ/`W��u�+�2�#<�ۑ�-���Z�|_��'��+j��o�GG�;�fƍIl��K8���Ś���?x�M-��G����0#�]��0��l%U�����f�����u~���Z���W����2�!�8}�;)��"n���	>{��V'T��`i�O�'.������P��7��;R�+`V�Ud��MƱR O`�i���?s��w8my��y�k Lw�O1�DGB�K�W�mOD咭��=��"�@� ����Jc�����]p.ȃ���e�&#\�T�g����0aF�_L����0<g醕Pz�ϪP�|�A��>���YY?��<r���/X�M�m%�S�R��\��pq���n=(�#�Ӝ�������OT_�`5�3� �����n�i%�o��މ2u,�p�ӬR2sS3N�]���ʭ�`��,������� ������N�46����3��Y�(h����)i����W��F�-Y��Y�3��Zlt�	�4���sZ�G.�ͳ����}�#=��ȿ��v�@`*�� 4$�ɮ��#<1�./�{��b�+�\(p�,s�R5���|�_6��{X�A�
�(���W�5"��f}�
�|�}��z,R~z�~�>7�	�	�s�lH��5�Z�i� ��}6F��)��y�F�IBX�4|���:L�.7�I4ǈ�pIR�H�P0V;j��vu�/A���sGW�5Knzs2x��N�I7�.�s��L)����$�gC����<�`ܫ�N�	Y�n
�M&�[û�7w�$G�*ȩ��Y�����{~΄sj�n���X��{�v*Pl������㱳O�.n�Πg���5Y�5�Uܱ��qw�r��ia�"�юd���
����1����79�\�e���H.�.9e�_�oEq|=�Pt�/6~X��"��;fk���Г���	"����Q�s�+��=��'KnFtz��W�p{���2�;K~\��J%���j$(���m%�,Ӡ-��:����q�-qμeD���{?*�g���ѵ���l(�\��z���G��!Lx�w�ob��]ɺ�9��And}������̤E{'�Vb;,���(��������r��҈>�;�I����Ү�k㗋.��L'���V�pI��Ga�����z� Y��M38�����^K��|+wڧ�[:tHvƈF�L}s�����F�ōHБ��D�̹�g���i-���)P��ɰ�{���:�1Qf`��_��lӓ&R��>fG鐁��f�U���LP�fs
�q|���czN��#����^k�ѕ�q����;�盧C��8a��+^�h��
��(zb���>-��=�+�=�9d�@�a#iyouo��U��ZM��w��D���#��6��G����$��s٫m5ۢ�Wb���j�[�%�(˩'��L�����R�ڸ���[т�4
'ϥI �#E!��Yow�p��`}̐��}��M��'*�j���u�.MD4B����h�o>�A2�m���D�����ح6��W���Jz��r9�A|qH��j5捻�<�?P���E����ıjoH�3�^�>.ln-��I_@#ve=�Y�V���=?���p��#<��#�1��%�W	i3EU���8H���M�����D�G)0,����8�i�T2�K��f��3�U��~�� )��vs�a@ù����y��]��:bxD�I�U��x�����0��B�i�p�YI4����䖔��vl�5A��噿,� A�ڗ��Ʒ>�M��<���g&t��F�4������06<��`L�a�?`�,Љq��'��|yP9N�q0'�
���D̈́o4��8gA����Y���L:e�@��0%��J���'����!�h�!��}?ߣ��`�c���,��� ��a�K���K�,coZ�\��۞:4�L�E���-��*��z���6���eeoI���4�f�̸!z���8vˇj���Ӕ^��5�h�?ҵ&L����މ�a�����rjB�;հ��T);��'���T7���"z�O\� ����*i9�r�O�.힌���ʊ�����	�2�`?���&Qt�VO��,�ry6DU���~�?��uQ���N^����'��5%y�\]�MCh#�vJ'�|��"Q�q��3-��Fw��dݙ���=�6�:w'/43�2�{0KȠ�W"%�GϲD�/U�مj�V�'QB&�q���|m�u�#`��r��$?"H]QY�_X��U�nv@'�c���bVt`"WMj�������}\�3<`d4¤�>Cģ��c�-r4�R�[1��3A��o�ĸ�"G;�k���y��Ñ���K�-�&����\m��D��U����=Oз�o��°��Ç�A*uW�I���)�vˌw��P�C����[����9��ns 6{�" P#ucf���	8���2�4yP����@�����Wf�1 J�|��^�D�b���}�����F'�D�!����p�;�wJ�W ��"�I�g�Gi�j�O���qaG�/��ύJ�!�*�DVN@�� v��k,��i�	�\��n�A�kB|ﺐsS�Q<c�E���, �9ע�m�;	]�WoU8Hi��\f�b���T68�9h����f/ڝui�S3�tv)��b6��,�5�Py����^��+�rC����_�K;���wwF�Y�k�W�Ά� rbG��L˺�Sc�J�Ɲ 0���",4��1�jQ��~У��.G+[���	x�w��D����sX�7ISG�r�k��+��'���2��6���f�E�ju��l�4�$�b�v~닩OH�W�������e���S��- �@?h؊���Szc�W�ۋ��X�t�a͓�@���Ѓц.5öMQ]���$�yIP�h>G���hu�H�>����wI�p���,9��N��Xjim8����� �y�X�Ϧ.-�E͏Pfh���S��a��ս�����h�p�b�(J�����6>lIH���[u1��/5Lmf)������������@�&f��:��C}}|�%M��C�<U(���)PW���='UK��������f�{Iy(���l�|`q�D)>���(ԯ��`M-��Px˓E�%�zb����9����J��b����e�m�4�(���-P�od\�A�n��A��Q��ل�N1ɩ��3��+�+ɽa�U�����o��l�'�p-�闠/�����'^h�g��w��^u�O	��������ƞ)�q���qf"$�y-9 �4�\��J�ip��48dZk�4�@=�n,������Nze��B�28+M�����4;���z�n�B��ʳ����1��_?����ߨ�q��.�ʧd���ʙ���9$�ߺ(g�'���oX$3ky�Em�j�7��"�N�D�]C�u����B�������6e����FΨ��k,�聾� �Z�l�xm%VW�Ld��]�gH1�	��e9�d+DB43��<n�K�8�D��!%�{�{�����Ϳ���D���!6��ʽ���T��DT��L��|�aǯ,�m�f�S)؟S�����-q��V���ec{�\UER�`2��"�Z���{#�z��X���#޷_ \QS�掲��-vݰ��1o&De	U����������<��������g�/Y."���4Y�n9�0��2�Ǣ5! ��=�@AN�� �>6v��3��D��7BS�%רP��d��i��[�*iMW���F����.Q�^��4B�@���1/��}@�w�QmV�"	���������r���2zp8ِ̞�Y���H8y�*��%�;2��f��"�U�/H�@��-�ܛ�j�`kӽӞ�E:�\��	$��}Y��LM7,�2u.���V��!��2�
+�[�oU�����؈�4��4q ��@\�$��n9	��)tp��i�5��"L��"-+6�ڇ[|�����ۦd�8��=�+3d�L_�'b@=�]�Y���\gR���j=��� :zo�§x���a=�32��oP���i���%����wG�pv�t�[{g�տ3_�ֵB��g���ة[�cpi�Hۋ�o-g�
�P���J�������9l<���~��3���m�=���w��VЛF)�m:�͞����4��V�ߔ�l����q~��;���[ĵbeƘW�V2N�:"Y��\��ְm��G��qga�H�7֥E���a!��`*�}�1�������ې��y}�*�l]/��KN�u��y�S��K�,h����+ ���a,�x]ҩd�"3DHd�$L�	k�
1W�#CAq��Ck��ڈ�8��3�L�W��\O"�A�6�&'�����w�Ě�?9ٝN�������g���H�jT�4��*��!A'J��YE��?`�n�><�ے��3�1JT[�i��b��Y?�i<��Sp�bf�9�[]�������|AZs[�C�GiZ��-��i�Һ�B�3!˓wc��]<�v[kZV�(����"�^t_aQ��*�l�$#Qɗನw�u{I5�'o���k,V�f��X���H�`>�pT�ft���01h��O�	dH��� zD��C-��I��"7,�:/���:+<��Rr�YH6[ew��)�D�n�2�Z�!�}�r���Ht�f���m����� #?�:J u��*V���;{�L�>���|�:��2�;JU�u,�����L�~dr�<���3������G��;H��� �ti0 7�\��2D��>4��j:~_8q�>^>�O��3U�V�j��M �f�q�0w��$�mz��nls�ߖ�DE��9���{K�]�1�����|�Q7X�:�;��>���(~-���޴�I`3�pC���(���dr�5��Se6��^:��W��('IPş��8X���|��|Z��iP�7u��me	"�%���yltM��yؐ��k�ߧ�Q��c��$�YN>��a�E'��>�R1��Y@�[�a�ʅZ*J����-�E��}I��~1U��C>ΰp�Ҫ�>l.6���V�{�Z`�w1ݢ|:a����|�"K�ĸ�IJ0���ˑD��$O:3�BB
���1,����K�a��t�u]<���2ݝ�O����fi����ѳ���ikV5�:��'&�yJ!��¤1b&�慖�$*]�O�mX�� ��E{��[m�:�A�"�$�(?,����f�j����1Q2�6Π{y`���̮�����^� J�㿭� ����[��0)=�-RL���V-��։�,^�S!�L���	.���Dt!��.�<�EA@�8Ou?(���ι:<0PЀ��S���w�l�NV����b��6}�B9���A	 ��O! ���3��i����J�4�.]���{1��^4]i�J�8e_R&���9�=K�V�S��/�ìz�"r�&:*��\�����e��C���#�&��ď��m~>^��y/Bi]�m��G�wQAޚr�L�"���M�e���a8�,���@��si�^�PЕ�o��;sc[Z�D��"g#���`�8�������R&��=z!HOsd��-� ���(�B]��r�^������������,R,`.��ߖ�f��!8e���]��n�5�]�c�\��Q�n(ws�VJ�h
`���������2\�f3�,���l�Z�B��	���U�
x�+�?�]�G}�`�p 2H^U�-����'3�,��ݥ\���~�q /���"9����	GFv[*�]��@����ۏ�8!x2�5���Y5p[��_F$��~ـ!I�0��_w�������j|����ҵ�T��{^&�ľ�o�83�񈻆/�@y�_N�v�����O���gl�~;Iҿ��ThH�е��|�OQ�ے�T��"���g�!tO��X{	y�=��~���x����d�DlB�uĴaL��iX����F��'	@::r�q=�N���2���J9�Χ����D���Ŏ��i�sl��rD�id"�`�1�ȓ�[h�����~�.�=�d����'�PǱ'[���=Tۊ���#�8�8g�Fd�k�Oq�-��4��S9΋���,��Q�=x�'���ɨ���B�������3�nOk���V��ײ�j����%��*��u�7������">��ya�ᡬ��Ķ�O�s�w���$���
�lV�a�O>Z���"yvR{$�#���g��Mi��߲x��. �����C�e��6h�1�R4+�Y�;��"�K�F��r
n�}�I;o1w�E�����c�g@��Sm�Bipj���-H���\���z�Tihl�좇�|w�
M�ga)��+r��l���[p�m.E�\;���n34i�����֜�б/�itj[�Z�ь�o^��O*�d[�;E���Oa)�(T�x|�Ƙ����cJ��&B.#B�E��jk>|&����h�>}�l���ݰV��l���~h�J�����)����Ú1�͋������Zt�����/�b�X�$��1v&���;����#z 4�KB��$I�3�L����N>_\W�o�̩ޞ>Ћ���3��t�И(d)6��`��x��ɩԴ���xq�����϶� �:�l:3)�J�N�i���~U,��N5B+�]���3�}(|�6pwy�����c�,4_=$��L�a��V02��Q4z�=�vh�1X���:2��E��s�r����K��Zn�B�Gm�(�uC=�1L�i�K���!��?WK�9�����#����.%Ԙ���	}���N�l^:����$����<_��}�Rh^��y �7u�\_�!����[:|C1�3�D����^��=��j�륍x�8j
���A�F�F��!�x��!�vD���Z+z⇽�e�H��*�\O8���O��6��{õ_�'�T�oz,l|=�UW�N���\F�Q�F��ŗ��Ƒ���-��!�4N��r`8����!LJ��*+����.��9q>=��h��EBΟχFe_���������Zg�w��������=�����B��T�t�h5�tM{����L�$���������I|EF��.�I�p�Y�x9U:���Y^^���t�g��+d�"x��N��9���#�$�&����u�D�ͳ�'>�s��(�=w�$�5q�L�����۱�s�,���w/.j$���9�9�+���4ަ��qW�M�e^��ȶ⤪E {���r.���r�`6�HaY���*j��V?H.wD4^����c��&б	@R���d���dn���'��O�F�`�@�66m��IO�.�>�ȩ�N���Ǥ��܎Z�8O;����842���1�?W���8��y0}���fi��"�<��x6iWK��x����Bh,�K��Ez�����O�F��	���m[~m�I���s�\�i4 �  ��`<#�x�NM��'�F�X�w��I-w���`Jj�Px����ˮ�"����C}E�G�����G�fV�o)Y�,ih@l�w���̏����L��
��	_ũԱ�*;"NN�w-B�f��F�w{%`4�&�X�B��4�hJ��F*��C����N�I���h3��gP�P�oޟ�&����H-�/���-���E�_:ϫl�.�����T|��G�]�Lt'�J<�}��ʞN��#�	Qai��x��1��O��)�fvf*�;T��%bl<��r������`YU�����g��(b�X��8q"j+ƅ�9NOk��O�L/{Tc l����������� -���3��^��M����HԠi@�>��"�ܒ �ށ����$Q�,���=��$��O�>�a�ŉ���)-r©��P���Ҟ�I�Y,�+�7\-���
p�PA����я�Vޯ���%$��Hh�pV���X�Ϡ���']v?lt?�7<�?EN�m�o#��Zf����(b�[�$x�������=g#
-����N��,��2�֭��%�SdZ�>Y��.��dg>v���z��C�r�(�����C)���MZ)�v*s�����������FI#j�=nM�D��i�J�۞���NZ��E,�u�d�q�̓=�����JM�%��iA�c۸��w�E�����I|�C��4R.�:	�����X/��Y��[�����_wO��HKzy�m�0��e�?�����ڤ��e�#��e���F
k$���<`JL"��-*��y\��4��8?�gF�@Rఏ3�Sy�F'��B�'�Y`c�Nn��Jb���*� ���	xG�GM�C�NN�Ƃ>R*Y����Nw�p$�i�ʴ��cǻ>����u��ю#:r6�t�c?a�\ƌq�c�L|pUK�.T	���۟�]6�	hq��x'��'_~C5׫��V.�$Bf���!�[c�?Y�W�~q=�=���;���.+ܚ�m��A�C~�N�*�p�A%Ÿ3VY� �t�p���/�ެ�Ԫ�ƃ�1�bN�[���S�=b��W΂��T��HP�?�bh�|!�4���S:��"�d��H�ya�W?�j˺ ^.P�w���GAQH������U]/+�
�tж̀��d�|��}�����D���>�P�[�#���P��x!�sڤ\�&�]����F�Uk+S9���l����<��{�1+~=V�d.Lv��aZGM�K|G!i���N�s�&
��0�=����)�n@]�0&��<S�4a*L�6�z:�b�
����k��~C7����-SP3W'��̎p�Y��Ŝ}&��T��LB٥���,U������P'��BW�"8�je7���E 1�9X�7 �+��ͺ�:����1�^1�<)ڷS��X--R���&�=]f��(�g�^]��m0��|`�����B	��^CMH��]:ԄB��:/�q�ڟ��wt8�_���J�K\s�D���@�ǎ5�i�l��h]/��RA��9�7���7K#5�I���@m��;[2��
{�L�l�w�2t�wCMp�+�%�o�[�	��7[Ԁ恇n�W_��%s1�����2�C ͟���*��j�9�?��XE����k?1���a�$_n���Bb(���Q�6{�<�ԢN�j��-l���3,�Saip>��k�*��ǔ�W�9�i#�UJł�C�z����P(Pʔ�-L�+�*�o9��)_x8[�'$�K�y�����؏�V,�X���|u�zE7<Ε����5��G�nۉe�s܏�	�*�w����Su��HW^�8I(y��
����6;����{;Kà_5���Ϻ�����'%~��_��'� �e���]c��
�E�x�ISX��* $bΕxz)�������$�:ՌuX	�N{8�ԝ���愐/�^��!�Xe���cI0C�o�}��7+f㫦�Sa4�dc���S)6%%�!~�p�Q�n��o��H����r��];�o��Z��#��Q�J�M��3�6��B���o��r��"*�e��A|�}r*5`��\#R\Qbv�����`dHB0��%�*B/>V�c���
����O��p�(������X�S�g��O6h&�k�ʕi�dj-�:����[l�=V��Q�nsO#��c�WI�.�U[g�K�x����{�+�x�y�*��.]"�X�.�s��LǇ���y���Q�rt���O4m�X�<��p���+����%=V��L��i ����͂�B`��&_E�����e!vm	מ�Sd�l��O}S��Y:!{Ր~�� x5l bM>��3S� ڃ|C��\���u�D#�r�f�Iu*���O��_F���3���5z�[��n��]���� �ق�J�4��^Av:.N�Ҙm�}�Mqa���.p]��E��q�]?�g���d#�a�oH%IKLZ:��ƕ*��	YT��1�5����p�߇�I+cA���Ɉ?��&iŏ�/qtqsX�^�P�c�~�Ml�(�����2Nyt�XD�w��|�(�D �c���f���0�~)��U�å��$�w�v�u��a��yV����A�S���#�c��3|8�g�oj���	���+�bK�T>wi�.zwDv��.Z�ˀƍo	�?J��-��Yj�m>�^�1mCuP��g4�$Wz���}�Ff�!P<z�9��+�m���m2n�[5�4屓��W?j��e�s�1�����^�
c�/.i\��r8��U�h,/w�Җ�{�~�ԭ�h,p���\���5Bw/�Cx��������Q*�׏ӂ�,��3+D�lL��9��3*��z@R�Շ�7h2T��3h!5�&�#HvH�\$����/�T|���������������;;��{%u���vN��uWS^�,�.��>Q�n?}�5�i@@�kw@\C�'Hr���]�[�ej��Qyʰw��W�3w�p7��3��&���W��i�}�#Bq�����(� ɓ�U���<Xt��'�"RF8��[�h��,�0�~]{V8^Ay_QO�cA���m7�e�}y!mt�ɛ<d���0��O*`�?f�VJ�q"sf%R�^�=�+b/��q]U��ט�\pB��SU��L<4��޼T���ۇfK%�m�U�bt5 ��yw�lG?a�Ǩ �$����
i��>@�/�/c �'�J[:��<�%ӵ,��H������r4Tys�q�P�_7Zi\.�O�\;H���%�rDdT j�!y�xX-  ۙĨ�����J
j"�Y���������$�bm����ɡ�r�k�\/um{0Z�9���x�>���l9�2w�������lG�,�b}��R�;}0���^����Kا�w/��1���S�BI�F�8C��[�������6�� ���f�t|�� �rEd�7���E��vf40�&�ou-�{c��zj&�����<N�Cu��z�akr�,�6"s��jOt�4hD�hodi�.�v�@��N���cs��m�#�.�8d��l�!���)�S9$ڞ*)�}�B�������(�Ck5[�`F:'{��H�&���2��P�6m�*ͬ�%�+#d�F4.�[���dR�k٪��n]\zȮ~?4Q7�����m������b�b*�r�:Ռ�I�P�}-I}��)'#s>/�Ӹ9�$���R�h�.�!�(}[�5*�����`KZ<1�ѩ֣Lr_4��fQ�Z�k1I.�RF�'��y6�t�ܘ�f�>
��JS1�ժq��4j��()#���R"�K�N��\�E���M*�ܹ��(�I��*�Y-@Ҳ�њDh�G�G�u�Mػ{�kKw���E�<Un�#�ϣ6��K���IW��x�{�����<p�!�t���	p<p��`?H6+w��G��6��e���-#{��Н�����ǻ?�=^�m�����/�I9�I�j� �Z��$E�&��W#o'k�1;�A�Y�.A���!��ϫKb���T��%�Aj` ���f4��H�V�"���5�|O0Ԫ�H����R@9�xǎ�6����ќ�����4ˡD	a̪�ѻnN&��e�?���q&���&�}�+:�޽��;�i>~R6����"7���0���^�e�E5�� |��a��6 c���#��2��B��z\ka�TOsM�G�5[i�:�TP�Ӫ(mh���_�%�F��D�	�+gy��a󅠳����u�6�/���\��+����~x���-�I�|�s�~�hQ�����r���-�h���}�u���7��Y�� �eC9(@ t�Ӊɲ=w~L�_��A��61��mK�u^N�f�rVA��e�}~eаs�&��ґ�5)T{�tӣ5(���F�l�8�w����,wD����� ł? NW�f��Go���?�5%��l���H�����i�%�S7?������b���P�41�p���P�)׸�M���^���*&���o�)n��^n��t����T�y֊ў J��q�֧~��#����A?��f�唷u�#���ϊ^���5}��{�9+0����XOЖ
�Q~��e[�@�x�NE��B+̂����o��F�ܾW�i?\�GPՏ�,�*"#�Q���V�@�5���dez�c��w�[���.A3}�@C�"���C�n��5���>���w����S�*�[�p���yHI�T����\[��m���X���ȯE�������5ޙ�߶`�������B�?���C��9g�`$I-��P�0�m?�;�8l�d��>B�d�q�N����/1��h� &n�¯��K�����i��eOX�3��>�^���Y/յ�r�{���͜[U�^Wb�K.rg�1��N�X'�&E,?P�@��|�+�)l�M�)r�X�^$�w�p�_�7~s����2��Ǒx�`����y�.�����癖�?�R�|�߽��U!� e��
�TY����"Ts@������wx��`-�d����7���\��--z��a<IR3]ly|%�/�e�]d>�c��).��Ϣ((����f�{�W`��h�XՉ�s��,�%9���}���й�4�bKL[���"����~�p?!BTeI*Z�h==��m��B�o��@@�񮷭l��V�w����uy�an��ʊ����؅�l�B�U�>�+7"���3�.�-��[k����
� �V�[+�yx��xZY37T���lA+J0[o(�w2\Z) A^�1M���pܖ� ��AuN�W�* ��2)�Y<f@̐�7|2���ۜYe̪����v{��@I�O��''�����OC��f-!@[����4K*Q��m@�1�o	�igͪ~�|:�5�l��l�ĝV����s8����*"����%�o��
y�|�����(Wu�!K����f#~�Ġ��#!:�\��xS��y����p��k���O�~��~����$ͮ�	~�O-�����|�W�K���h6�ϔ��L�NC�Et�3Wm繥R�y	o}0�ڣ+�����S�}} �����*��z���xN��=
�
���Ö�F��B�,Qb���ߔ�$��,������W�d���:a���;a��&T]��QI}g���z����|���"���g�RT�8Rv�-��<]dz	S�Y�՝��������Q0#=`��J���"�����ɴM_�ׁJ�'&�P��c�"��t䬿eLϓ�8C}� ��g���7�j]v��Kp���U7e8%/���v�QeOy��q2b�F�e�p~�p�����vD�
M�R�;�Y��tИ��)�)7�����1��;�`��{��i�6�̺���L�䏎�>�L�r����K��.r9a���*����� }-)��ؓ�M2R�YE���iI���%��Bdr������0����ЊZ�-����`M�-��"���k��[(�
�j�-��c��WO!�ot���d�l�Lf��2���t�cϴ�3����q=�P�bQ�E�'�ܦ�|ZX�}J,�`����2Q��!i���?#�1a�� �R^%A�O��0��H��d�v i2�e�@�PN�����M�gp��S��:bj��E�&䧛#A�	�	$���+�II��.�D9���Y�˟��ʒk��u���_ϡ�;l o�_���)ը<6� ����݅�~��r˭�oFY&��76=�_V����-"�d�2�H�PO�B���]��>����]\6^���~쨡'�Ӡ��E��SD��`�����J'�;��.�[�"���ࡌN���'9�{�܅鲐$&WGH��\��8�F"F.��m�!�P��� �y�{	��`�)W���Ynyi����}0��׍�Ȟ�֨|o'o瓳}x�c�[�ȩ��/�pE����M�_ûW�6�M1���Ğ���	N�4S���Fbr�e�]flr�ߩD�^y�-�p�@���9��:�Mp��g.�<�gP���;C���Y�`?��r�%S��r-���9H���D����]�'���t,��PmX6,��~E�Tu�A�朎����C�O��scH`�V��ԁ�P<T�h�1q`E��I�E("\pvm�iye z����O\=�#J'�!��)�]9�u�� �x�esM��ϓWm��^+��5�[��"�S�X���">�4Q:�����1����)�Bǫ 	>i]�=��1}�����]]̋�ɴ�/���H-���C( ���0�̩��� Hk�o�$�:W=!�b�%�� O�?q:"��o97F�|5ۯ�b�VV��#���^�V����7�� Bj$��&�������q��a�X��R8A/�CR�t|;~]a��o|$�Qv6�B!������
�;�E�^WU<�ӳ7rI�YK�/n��BǠ\c�I���t����W	�K� a�EEŢ��c8�JLQ��?��߂,�۪\L�9;��U���0��qD&M/��3��k���G�4v+�-*�D���+"��q*>D�D\�Y�+�be�"o�-�sO7py�Hq����!yv��e�0?J-�T�����F�v"�-�ݫ9�Y%Cn��y�l����T��e� ��v�(�
i���羅�w��t�#\Fʬ�}�}��B።`G��B�E��0/D��%�`@p	֨�b^�zF�W��y����nș�1�WH8`����/X�<
�N�vڼ���cWNa�2�(�
I�v1w�^w���a����)�S�XG: ���$Ϊ�2��=�)]���tೱ�>�����Pw��c�gN��Ʀ���`/p�	A��o��Pq�CU���}[�D	<7���h�T!�AT��p?�������'P�ڙ�'í� ���NA�i��8���Sƈ��]&!φ�����6�K�Ps�0J��c���H+��ɑ��ױ�z�Ϫ�h�0�x�L��1���dc�Թ��x;����f$���UbdC�ݭ;�Rl�i��vл�}����oz'/���;�tPN������6c�~!���^���ӗG��P��擪�W�U������ry�&+�a�ɒ|4�`ХP���'����=��BK���g*��u��[�OA{6�e@�j��_� :~n`�ÇR�Z�#
*H)�"� �C=/�Щ�^q�A��S�~�V���{�&���=�w�!�
�����9H��x�sBٟ݇�����T+��X	ߞ���>o��`�YD=Osj�-J�������e������;(8�M$�%�k�o-�2�fZ���2����}P�0sIK�&��ہ��gT�9��Anm`����K~�2��J��:cU���A�xX�-X�����d���g�,�"`�j���|�r��8��cG�����h�R��'}����
$�d�X�����W���n��u���v|X�W�p�5`nwω�5*\33��Z��<���S��u �=0ʜL��*x��uj#���!�"1jh&���h�go맿���X��}q�0�v��Qv�������7��9Y�%���ӎô�6fȉa%dŪGzI��X�w��l�&r�_�kY]0B��Q������1�a �FV�&��O6z�/;*���l�48s����GTç^��'y���V��͢~����_1\�MJ�S,h��RHUt��0�q�dC�W9��B�_��;�	.k��sU[���׽b]�B�Р�����<@��؎7@���
��+q�<c�8��&�H��"� m�6�<+^\�>��$��X<�n���� ��mǁ�H����q�f�Nh4`X��䬑�L!���e����\���Ɲ%�5�%~#��l�<��l�(}���'�(����ap[��0���:���������
�z�#��0��q+��h�aʋ���KAf�<�d#�ڵ�W������--�/Ɉ"�p���h�A��xԁ�������u�@o^߸��[q�m~��ν�<z��Z��z�or:� A(�s�,��^����"E7����l�T���v�y�;��#��9xE�����l����r�%�Y��
y������	���wy�|�v��^�>���V�����ʕ�o���oby�yh����A�_& �.�]�R��]Ns�9�N����K[臐�(��Q+�Oܔ��>qb��<y9��Zo��<=/�v��'A��\�� 3�by� BX+on������G��@��.�Q��Z1X�n��cl�F�N��ٸ��n����Lʦ4Ҕ+�\�*��$0g�,2�݅�
5�ǝMK�4��"�.��?���j_ZeW�#�)��v�{ɄB#���2�H�J�g�ER��#��-�^�K�tb�jA<bb�l|�U�:��������0hM�whK�ŤR��fbLw��w�ג�Ң/��s1'�Gڱ�����k�,��|��Bn�c#���$:�l�1����.?���ʊ��b������$Xa��s�kx5X��6f\~��}��PA�C�W8����<z'!�k�__M?��@�s�@V�2�d�f[��ɥuJ�{��C`���X.�Y��<^
%bz��\*��_	nY�˵��K>+��zP���ԩ�M�.���X9sXT܇"ʘ�AE�>�����WX�'3��Fsz�/�fVK�SP^E����O��x�-� ��������a��t|����i;�Z�~���z�jqk���+���
[1�r��56߫�M6���AF%g�@U�����yяa��PAtx�w®\�	��\A�o���5�g���!����D 3Ł����ѿ��b/TP;߀�+Ȧ˷]��F�<X�$�U��!q=�1z���D׿��1�����V9B<�m"��IAXN��V�]{۫�ڵ���vaڲ��k4��zEi�A���jdγ
�3�~a3����O� �-�4��=��#�ih	+e��Q�!��A�Ϭ�g�Dv?a��o�=���D�-�>Jc���}mr��ϻ�	Rn����C�&�k�:������4��`Kw�K}�~]<;����	�0Pid��󯝳��mxc�5/Ù�Bk2./ݝ~tJ1���߂�����`R̸l�>u�4LY�G\�0��`��\:�p�'���4C^D5�h
(x�;U��Y��N�)t��ߝ�,�b���gux(^��GӐ�gmܪ��~�g��ٛ�k���~�?�5P=]��x��/s��fZ�଎��%�NF�,��Ϭ#l��i6�Yu��������ݢ�@e8O����I�����>�G8��°Ҙ�:�U�o����Z$�8�l�	�A+*�gd,��)�x��T���Ō��;#\�$H���X��'?x���rr/�PC$�F劂a���؆�@�8P�:�vY}X�ɁYW.�^��3`0�Ҁ��JO^�3/_4g�8|�q��W��z���Pz*�E��Xl?�G�f�K� v8�v�1�/y��"0<>���;.�Yꎱ�G�j���,��{�|I�}=��\���ԭE]�&8�l�0C-��Q������l�����-����L.�&8�W���Rf��anBGS��a��0��2����88��v��v�.˼�H�����v�.�g�h +KQ�@!��YD��n4˧>�M�
CYQu]Z<v�*��ҧnva��y���L�Y�i ƨ��o��M�ȕ�JKHZM0�����)�,(;�8�6�����md"+�M�45�(�k��b���J=ň8�q�����""ؓ>���vմG¦����npI�n0{=c���U�7*d(�����H�e��Z���ŏ:	OM�
�YQ�3W�H�=�=\���]8��[9�qt+Sc��YZF+��5�Wm��I\Z��Iݮ�(��^Z[Ȓ���ѣn�<��ؽ..�>-����d�J{��"�F<�*����ʅ�n1�k�1�ŕE��QF��*��dZ`ĥ�~{�u��D�PRs7V	썫Q[�i�����5�7���]�B�~�z����f8k�8]H/��_�b���_�&���� �ja;0�~����Φ�Sk=U��Xfܔ"��şM���V,4[�L�M7����~�T�)��v/E��ў=.q�n��b�BNL ���1؛��i���d�5	�t���S���a��K4�8�4�B���t���(�Gf��Y�|r�j�֍=ų����$s�H����j�h� .�9��Z7&���CkXO���I��B0�����v,B����ݢʿm��l��>�s���W�D�؇!��C���y.VN��
�.�N��������dn���7��oI�]G���T@a�m�B:��!��6����M-t�Q�R0��X�4�f������N����?�O�sx�&6�g��A]X�^*��?��>Z�a��ȴ��&;�أ~���P5�e�ʻ���{�����W"���{�x?@���n4�:�Ѡ�W�s�,a���	�^M��.� ��{2�Q��h��X��\̷u�|Q��z�m-4hpĭ�gԂcI �{�.vٵXf�a豎������;Ċ�iKJ��0'���`��|�&��ɧwF�{b0�*�b����0��T6�^���"�����`�{S��*Ү�^w�\3ʗC<�F\�R�0� ⍵�	X���r��H�j�Y0&2���Cc$�U���|��#��VcQX��~p�U��Tl;h�b��i!K�4���ː�jb��������\A�oT���#�Ѹ��RD���M>u)���
�r�0N�v��b�Q�X���Y���A���-���#7��3	�jU8{\6_C�א�r��7��l���B]��G�:����Μ#��<�L�_׋ :ߢ1����R>Q1!��f�%�T�a��}G���/U�4͛LMqJ�z> @۰�fӠ�2�Ė	��d�_;Ÿ;��XQQ�%F�:}���P֧[�|s��d��OK��0����*g.*��P�{z�׉o'_��l>�LQ=�9^Ҏ��M���s[�4��*@�4�%o����K������S$�j���O�@��=Xd��=�J<�C4��ǫUq=��i���,�5���۲�-E�G�y��_-l"۴�h#�8H�s*��1��^�6���l1�e���q�E�3æ�n���I!�W��@��ٯD��`g0Eg����ʶ�����8gQP����f���9���-���l����?	%xk�l4�w�-�+���&> >	�ˍY��������h��2�B}�OQa�'q��	L�6.i���ψ|D囘��z��ڸS`�s��6L��\˙V�z-{����}5��|)�Ϩ�"�*���4	V��d�^��C5��Ջ�N^���5�D-L��޴=h�A�orc:�]����saS��RFUV���,�=�s"���s�g{;��tM�M��wV｡���ßaH��[�$��id��<AvQY�
p���#�$ҋfBC�����{�|��jm�aWf{������e���`��)[k&Ϣgun�r�骽1%1ȿ�)o� �Su�&c���6��k�m�-T�5">8��j9-�Ś\�k�`ҕ��}HXd�'��8��w�3�F.
���fZ�[��
4�-k��)��%� 
0��r>��y\�'� �I�߈����5��&�,�^�R�C�d��3ƣ�~%5�~d��í��^�����=�%y}�c1"��/�G�&t\����Zeh��!_���K��$�X��9�!�sI�Zk����0��%p������n�����=�^4EP�
��z�Ҹ��B�k��cxJa�_4�t��է�w�=]����Pj�#*Wb�'��+5��i �� ����S�7��
�g�R�";F��q�Z�V�N
C��Q�h	u64�2K,���1$B7�J�
�1��`#�.肆q4I(�#�����S=����߮��׷BI���c`mL7k�!5 ��/�Gy_g�r�,��&��H}�\�8�ΙU+�_e(�a�b��"��	�]n�r���qwʜ���͌�^̝��Ҷ�ꨒۖu�9c#���ీ��ȍy�Z��gh��
���>����RcJ�P�=;��p�3���C��-�h���Wm�}�8O�ć%΀�Z�����cy�Ҕ<i�!���X<5�W֐Ft�J�fM�_��$�.�|ջ]B��i�������h؀V7 �n阇a��l%)�W'u��
�p�j��$���x�%e�d�5Љp�Zu-*T"8!���Ō�!�(�PP���0�U�;V,�y���OP�֏x��X+���  �NF���� {KM�"�z|���E�]
��֢r�1uJm�A$�M�9�d/Xe<A�$���P�qv�*�dD��^�@H�4`c�:�e����r�u��2+~�'+AG@9��$F0�q�5`ޥ_U�\"�t0�j+"�H܅�&6m`�0�YH"�r� ����4[�:
o��'u��a+�F5N��%B5�<��H]���J*�^լ��O	ጄ6�]�����{�G����6W��:�ky��b��A%�� �ԾCG���ŉ�$�P(ܸ߫�]Zt䑾9"J�h9;�����l;��WNN�}'��B����� ��>3mGl,#�0.Ľ)�Z*�/ܞѩr(�c8N���G���p��7^X^���̑>)Z�n�|���F%�,׿����HH0��>�Pˬ�y���*w����%�R��̛���k��P ���0l'z$'�JUD�.�<4f�y����%H'�13D����K��HK��4���"L�#$�7_5?��	�_�<[��jX�H���POF����=���qC�=����g��Z�^\*Sh�(�#ޣ�.\�:#�;ɛ	,Ñc��^�����w,�d���PO�s���	�q��ɼ��y tD�_I��.���E����F�GC��0hz�l\��s۵H�V��2/6�Еh7�`+;��h=x�ք�v}�/f�	+��J���I�hǁ�����P���
���nwd�w�lr������?�UE�KL�pT@?�|�t&Ϡ�^ˏ��&)A�{�zvk��)��b��Q�ǹ�^\����8������,U%Yo](jP�ZںCs6�b#:Ͼ���@+�{�����C,�N�`� ���V��Hr���\9@Fx�.�&�_�p,���bos]�'�.'6��^�]�]I1�?pMcP�)��ܢ��Ե����lc�)c�+\��.T��E؋ӭ:�?�n����l0��	��,���z(̇69�a�6N��
��8�\���M��]"X��� ��G��lGe��2�[}X�)����wD�f�0�d�mιr�������٨�Wy����8�P��Rd\�J�`����ƺaqxBr��єm�:�V|���v��8��v��	/��[�hH����*Ѧܼn�u{�=�8����J���RG�gU�a*X�|���K�a�o��k���u�"̀)��:��ƫ���x1sϏ�|~������_A��9?%dump�)�]��+����m:��k^�����>�)��H�m^]&��&~����s2��H�14���vob��9��Z�r�ܺrvXt��u��Q|�6�!�=� �賲$�ŏ�R�+$>q���1�G8�z�E��v�e_����e�I�`�k��1Ο�����7g<$�ܒ��F�D��"��y��U�g8LW���HO��	M�A��:�1GX�;��O�^=R�A��%�˻ w-=�8u�i�7n= ��1�[�$�[tZފ0����AE0-���yl1I&��D}�1��X�11���n�k�p'p�̣�m�8���HaR�2GCZ�xd�zF#pSY�v
ş\|J� ;a�/&能���m�%�g��<&����er�Ǎ9�RSDo9*�l9fdkS~L'2��}�v�w��/I�u�~�a�~�Z	,�G�LE�zt��x/:��i��p�ү�����'o	@����+����/*:�]�ΛU_���	Z��݊guL��o���/Ό�+�u��閛RK�k��G���� F����QdQ�J���uZ�C�[�Gz[ꨤR��!�6�9z�ݙĳ��܌,����A�$	(�;Ц�*�`�^���ֵ���+���y��H�UUGAF�݌!����X�@H/Z�A�?O�Wv�w��Β�$���C��x�P����<+.�"��<6}]�	�j�x�z��Bz-���'r�w�����Nu	Ҥ��v�|�3^Oh;��5YM��ۘ�m R,�_6!k B}��P��Yb�@���U}޻]n4G�TC�+�9I��0� mQ��ԯ|1��aw��4���`5����P�FV�i�h�Kcx���1�5�>m�����t���{�?��T
�5lH��n�53�hy���B���P~[�
j� �ڌ��X�tb|��/���v R,.�I���6���`� {��	z��E�Y��Ԣ)��2�)F'v[�#'ְM�b���Y��D�kH/�2�q-��4#�NƮ�M5u�7��[�	�~�(6���_�	�����'�T���WM���
��_� '`��7�-?A�K]N�n��խ��Q�e9H��۬qȻf�|�|�~�9��E��SB���ŋ؛Ӡ�UZ���rk:��d�0���_�n ���~�t�է;�^[����~V����\4�� Y.=Nrj��gx"�#N�q�5�Qg�@�-�����05@���-	@��&HՕ��6U�?/�f�9����(�����O96�o'��=�ܱ�6ّ�]�P�RwՂ_K�
7�Q��52�#����b�p{Z��_TD�o:7e��ךn�` �����P�Uz-bEg�M�K6(�j�8nc�ėsb36Z�ő�P���WM�P�'��S�"�*���P�F������	a�cd7�퓡��D~��.�����MtX�2{�k�'b�Ɖ��0�\o�bO�  g@��\���8N��������mX_m�LR#�Ow�&����,��\��<�x+h���޽ދ�����<޽%>�������8�8)�����j8ߌ�8��a^�	7���O
.EsL&��1��yk�o0w%��:���lY���[����2��������l��\��p���Dx��mAg��(���d����x
�Pj6�$հj�a����c��m��h���%�n��0��1��e���K�i������tcw#�]�O�Gۑ̻Q�;jZQ�T�S�Q�pƝ�z��I���|˿*�MH���| ��'�@��p#q��l��� w��vB@t�Cɽ	%�e�7��r
��\�k�I��b�cA�OA��8R��5A�]�9)
���w����d����%��M��N[��Y�m.�1uIQV^�	CNxI�o~(�� 2TD�:xҹY�L��4��ev�-lT�۞s����f�f\ g�&�>��3�=��\�Y[V �X�Kc	l@�>� �谎4��0=�������xw	N�.�'���D&���2���I��E|4"צ|�e+tX5c=��y\��p��ʮ�;���&��*w°���p�_"r�����l�oe#H�Q	��~���N"?������dA���-$�5��܀ ���-W#���)�K,'v���ČtJ��g�T�#���&,̰�)��DU�L��X��͊#C2�wKCD�ej�r�B�"��H� ­�Q��g�)&"Z�Vun��N�������D�h]:��p�Sǜ�ynIv����2o��^�9�P`\l}�z���g���M%ش��5��o�8�_��/�~P7�#�rSen)���p�uK�����(�-��?��q`8�,y������K
�d�`l�I�MF����>FZ9��	G��P�E��x���s!������n���a��sZ�G�QRR#wS�^E�9h�n��U���e1M�8�RZ�tkǋN�_/�l����7�p5�7%��&��=l�~����nتfA,(_Ƶ��%��N#�a�,;�W\�c��(��)�x��5|R],�C
�É��Q7D�p��J']�%�4�R�&�!��i�FK�'�������SاF�S�T�|�b�s�<������IQa�AJ��j�ݢ�+� �^&'�Ɓk ~@�.�)7���$�8*�l���t��>��'��I�`@>V��I+���vE�����;��e��7�;�&J$�(�@q�!�����ڟ�~�P�F�o�����7熟��^=��Qɬշ�5C�5��L���
�^�!i�<�+�˥̪��
�A���
4�0a��۴n?S+w�<�)���&�낐l
vV"�}�>�>ҟ���-�-�E�y��^��$=��b��d�?���,W)!���77@�=�8��CG^��Og@�T��!UO�I.D����#��\��u~P��h��I�I>r	4~��Ơx\;�<�R�9�./+�8��x�9�pھ�< ��0��f
<y��Y@O���3���ܗ�� hShǫ(e�V��1gp��47�z?|(�R�c��^�C#��-=��	o�L�tD�; ^�~�^6Q��~�H�T��n�g��_#��%��k�/3MJ�űZ���R�I=��Uv@�L�0���є�}��Ҁ�v���-���i3�#fUm���R����űH��迤}�;BF��A����@D<ȋs��E �IMA����{�O�z<}h��T����e����i(2�����We4v�%%���Q��e�ۺ�'е;�w!��S~�P���7+�>q�Z�����a����Ԥ/���g��)�1�v_�h�X�7� ��r^JZ�3��[�.#я��~ЍAȨ"(m��ˊ!��qb� ;��|7� 8�e`�bɈ���Hֺ�&��m�dn��SV\���0�
%����?�	��(")	������ah0�|Ó�g'Q��^�+oY$OS|�����'�t| .��V��x���c[�FY�*�U��}e�}̑���-�D�)#^$��z�˳�Չ��A�"N�B�b��Fв}M9�Ϩ�q_��:�������2�%���O�%�	���6���dk}�ն�F�#�3#��?��q� |�1v,|L\��sHs0�z�S�G��F�dp�C��<i���?�I�V����/Hު�&/�3C/�P�ݒ�9\�6�K�ug`˺h���Z�*�^p%5����G�M����Z�L��&��v{�g�,ϵ�D�����
ju�6X�R��H���J��TB�"#B�_�DH2Dò��}Dx�6�O�:��N�#��󖦦�C�Ꝋ�#:7���f��XvPƷ��5���W���!ᑹ+�GU��N��;hw��i�V�Ȟ����"f�ǘk��z���CcA#��&�K���Ke�Յ�\Xz��ü��eP.Rx�cX��&Q^��]j/Y�ͷb��<�n���X+:�w׵"j��y���c�MYx��.bR������x\@�*�Z��'B@zv/���t�x{�Í|dP�R�x��4J1����O�U���=�/K�	-��	�܌&��i���L�@�2
ub�������A�p���ƃ�ȳ���FYNi���" q��=�0�RV{�������R� �i����ia����vܠ�cM��B4w�*�+2i������Xh�9��`����[�UW��j7�[z�=[!�񧢉�w߻D��4����lz!�7��G,ە�>�U_�ˀ����_��N��yd��%lU��~/�\��0C�����c�]M�TA�*�W�R���!yC*��<�a���������t�G�b��2�*�0#gmCKӅK��7��J���(���l�rd��P��53-���&A0�ﵣ>'o���9���2L�rܗ ;��hW
���aM �0 p��������}Z>O7=�)Z��Ɩ��x���7��nl�ϫ��:?Ӽ_	���}XB�z��Y@OM����85cl+�G��h-��Y젔���}>ԡW�}����ro*�ZT�9�������]��]��B�d�9E����s%�p��x�5 ���L�NB��E�2�
�.M���Vk��Y(��u[c�a������&y��`{gr�>/��r��.���E7�>��/U����Ii�2�����"_���Q,M��O-��7帄ڝ���Y*:��;�Ω�u��Ӳ�m�g ���|t��%�k��TDߞ��P5^����5��[��٘�آm�ܐ���m�A���*9W`�WA�_c��u��K���`0=BO'R����̱?�b´J���sy�U5��Ol�~��c�a%�y�dܔ��X�b�l�yF�ۈ_{*�)CSz��!oZ'�k�[�䵺wS$��m]\��i����� ~4XlPs։� ��Ǩo}���(�@Xu�������#�������L���/u��RL����2�`>@�SD6���ź���1������Dջ ��F���E�OvͪFj�g$����ð���m�K��(���$�"���zL��Qĳ����)xG��U$�����1'��j1��d�����J�U ��w�a����4iu�lE��j�1�2�}�鯋��]��'�ޛq�UMnd�wl��p3ᇗ�q������X�qp����!�C�]�q�3�!VJW�n���ƶ��wN��>f�hMBɢ8�z��op����)�7NCA9T��p�k�t�V�eu'�v���.Ϋ|wMK�N*e!��1j�Iq�N�Hnp�$��k4�K��aGs=��9h�lw᪷�(����0B���pp���L��f��]��~�BRH�ݰskMT�q2���C�E$��:��
����U�����^��7����\G+� �tvp�#���N�ޙRr4#�.ƻr��F�&�vh�(�r0�� ���ATR�!+Aw�sJ_J�Xڏ0�g�w����q�m����|Bm�-H���7�"c/���� �I�༐>uj������!O���NS�,�ǝt�'h��:��6�{V�x�M���(�F`���
s����'��q�ty�K���4An"_g����
	x|�0�H"�IDgV7�kzh��n��S!g�܍(^Ke�D}�]̅*�������;h6��Wȍ�E��'����q����|R���>F0d��y��n�e2�jG|W�/h���F��z�<���!��/�ל��U���N�<3v̫$�������|8j�P�r:�弚��'%�n����Q=;�9dp���N2�[���N8��t�;�eSD<�;���E������\IxZ�h��B8ҕ�m{�������8*2� ��%�HD<�E*t���zp�m��J��xK��^�IR�mj�=auC�[�4��n�����\��c� #�H���ª��0����98[�Z�f�9ޤ	E��iO�4�㽮X�k�F/��Y+�(��Ux߈�R�g[w����"z�Y
��[���+T��A,��-(1�B�t�٪q���Q���̙�b�#�Vs"VC�����}|�����@d�eV��R�L��R']Sk
FX�h��u�Ƒ�m$;�57���e~u?)Tq��6G����p���@݈(��&���	�Z��x_\ȡII�}4�,�H�Dh	�y$���K��vdF��skK�!t'�(���ćЏ��Sc�<:L sƦǠ�%h���X8��t��$BT5�{X��7W\Ii����!t���F)w�΄��จ�.
�v����q��d�,�K��C��	Xjg���_��j@I M���'��
$��!�_c�Ts8�UgS�M�$��:��GyP�kV�Oa����ɬ�P!G.W��H��󪤚�����{��y�(0칎��<S��L�`��KGT�Ug��#3��V7�3�$�|�����4wt���T^+b�F�fh�$�h`����81v@ʣ�?`�)����p�*x�n�zN��B����c������'�̎�f(�'$|��,(�x�����pQ�LNW��� ����ۻ>Q�w�4�h>I�mK;�b]=����9I9y13���7T�����痢<��D���W���������D��ϯn�9	Q�0��m��﹯
��;T�yO@���G�]��dW������У�T>d�XVҲ���{�<����#��q�3��ʑ�B+"�GI�&,�B�Br����.U7}
l����F�*�C�U�ڵ]�>tN�W����J����H�Z-V�kk@Y��>`�����o��A`��W���܅$�fGH?�8}3x�/N�Z1ʣ�W��i��`���q�ï>sC*�/b�DvF�5k�$ˋ�lM�;��W�k_��?;�/�QCt7P��Qή��izC�Qa�t�u
�e<ʥ�碆�j�b>C}��i�
�㟂�Rо�H[�z�VVM��F�@%tY���vtَ�Li{<Z�j0�������<5��Z�����U�9�kv��a^��]��C��p�B_�"�Z<��AyJ���'�Xv�ݘ���NΟ��̦ޖp���(�'NH�d8X��I߷B����\�*S��z
�4��R�L7����OE��e{��N�c�Ir޷苼$P�d��&�e�Ϟ��&�3Ub kt�M�[Ը����p:,t��݂��%Ht4�����̗�R,�<��B6�����5�>�	�UH�$�����MX��+���d30�SLL�E|���'�6V�^���1�n2��l0#s}�1����W:����C���(���Fg#�̛��LX�]�$�ǹ�����ҟVjI ���֛�����m1(���[�u��Ѻ���E�nWW��k:c�]�y�{�7$�^��96]5�����h���qFa�����<6D�gz��U�,!�
��;sJ�M	-���<|��t,������$�FrKD �����z� �/OL]�l��[߄�sV�y���os�������1���?�	�;����Ҹ���!�ɩ�v% �n�5o.h9X��K�ˢ$���$�zC<���v�ށ��G{`�]j_����d-	]xX��1�VP�Նx֔Ϗ� %���S������Za�ш�H�7vt ����T��tD������p��T�]N�ۄB��	@7���.�Q(i�����pS��l{�V����	��և���y��YM��[�l���I��]�����Sv�-����+ʓ����r�3�v�m���=|�c``�(�;WY�0�w��R� �m�u%u��E����Hd�%�
���5,���pd�^���i�͓횣l"�\1�lp�!A�(7'6�Vh��`�"[�~�B��
�u��~=�>q=�k��|�	���[7t��V��iE^������.��-��D�4�=�����z�@g73�sN���;w�����c�=�����]<軹3��]΁�J2i� |��8q,�H�73��
� �� �®�)eB�����W
�Wa�f8F�C���юލJQ>��ZnLRE����z�5 SgG%>�6=��LVZ�{S@�́�³U�f�(7��KY�"�õ^U�3=�������E�r�~*�����_Ÿ��/��D]���)&�.��j#��Q�Î�D�aj��(l��~�yw�$/m��][\ӄ�s�2(��@D�$�ɒk�+��@%^�����HR��3�Ԑ�cc3_X�L�@��=+���S��d
�B	 ��:��[{��*O%��\c��P,6�$�eI�ŋ��[���M�@���ZLň�,�6��3\$��<�Y�k�� �#7�r43}ϓ����J��ՙv�൏���ל�;y_5����$
�+'ٛ{��ڰ����چ���T6�(my���>B�S��� ⯼�Б��F[W	���rJ^2Evˬ^����J����0CfIWϨ⮸�t4,�sJWf��P�@�jHb�6����	M���EnwH^zv!�����3g�җ�ړ%���'�?�/ag�fR�M���9�^Q��E[�����@Pp��7��E�t4Bjm�0�m������T�赅����������p:83�GTT���.��Vi���L��-�7���p�6���t4$�ߖ��}]I���̟�:ʖ��T,j��~����m=p�uPO�F�d���=���Jp'G+Ӳ�k/cKb�/��k�Xs�[
}�{0���ه�7P28Oꎀ$�����L_,�-m���"�P��1�{b3��qE�%u��q��sxlqtJW� y�R'����x��hD��e~	�I����5;u+o��
�Ğ0�g� �-⩖��4/OL�o�
:���������w�[����$C�'�@n�m)���'}�R*�D�h���܍�����|����9��MLEӉP�(������K���/� �}�ʉ�w��"�J%�*�3q'��.eB�-�_>t��?A�
���G�w��bЙ�o}�PZ*5k��϶��'*��"���D�n��5_P���1���V��ߞ�Ё���Ue�41�P�Ƹ�{v��l���8��t��;z�fG��d��#k< �ܹ�B�{�/��1~�\�תB�.�����x�z�"�a�M!L�m�)C���^&hXp̨��Q�!pV5r�+GSh�Ԫ��L ��<�e&�{��Ձ��b��g=>�sP�����{���*'�0��c�O��~r	�C8h�/8ȧ#,6wS�4V�����e�X/0ɫe�G��ԩ!�9�8�|j:3���'��9Y2����ៗK=�(gnF�����=V1���X��� ��FwY�I�u+U�w�=��s���2�Ty/Udɂ�Pl��11�*�G�{�]��?o{9/��}��U0����`\]d}0���;^���ł��n�$Y�z6���&FUl���E�R�$`�΁����@w�Ӗ	`�����|?%6�lo�ͧ41S��V.Z��̰k�/� �j���Dƻ�~�Md�����X����]�y{�/<��m��p���#�$3!����3��3�s�`��zܩ
�{��?�ʨՙ���=;2"R�f 3��5�Mt�R�/�*���OAν��<Ս"`Wv8�>Dm���~3[���.n0���'�I�D��sb�V��"�kz�f�u5]Flu���'\լ1���-]��I�\(�Y��8����%��[��ğ��̓�-�9�AV�8!dS4�0TS~�2
�����$Ў!:p�We���d��M�ܪn<�M%룟�l�Y�B�a��Oū�\�����ĝ4-�j `&�E���s�F����jB14�sd�m��N�iR�s��?�� ������i��S��|�ך�o���_��aI�+	/��\�/0���a���B0�~�# ؑ;۷� �q�Lc*A�OR3���1��ۯ��U��Q5��^A����跹�W,�:j�!C=q�u�\y(|��y*���1����jvS�6�bN�Z�|�.�����Y�޻��U��hɄ�2�y���Q�J�{`�Kb]y��`^�8��2���u q	i�t���	E�7��^�	�=��ᚉ�����bĆ�L�M9�`& '�!hRr��b�c���I��vx?0&��9x�!h�b��5�z�D0S��0�Z��vm�w�9�15�'��
�^��e�V&6�๲7�Ɩg�<�x�?���cz���Uຕ�*�ORLD��xɫ��k#�'ަO��R�"����C,����wb=g�S�Q6�0��P���g�"�ZH�����vx��mXW5m�.-�ˉD����4�i���(ك�?�W"N�{(sg>�&����w�K�Ι�c�e��@�ЁH���kW�3xU�4�}s�Ļ�3a�>����������i0�o��~s�DD�w�,B��Ǽ$A�@�M�X0��QYH���g�r$�wI�T{��V{���KaיeZ�`�B���_�|���Ab�j�Ԓ-��N\�i�d������+4,X
�"W�s_�����kd�b0��o��h7V��Lů��Xc��*z�l��{U��F�b��A`9/En��l84¹)/�{��d����|F��H�]�g�e� {Ϊ��;�x�^xNe=k*�"G(r��ZV+.��)��Hk���׀H�e��R�O��'��,��t���dc��9�uR�dCi���F���B1m��pp~�?�s��mU����?��EQ�."9����Nd5�[�
��i��=DBq�^mU_��0T�$�5���$NxF�F�&�^�p�ֆ�s;���3ww�Y���4���I�t�c8D����ԀPQI*��7���5���*�k�y�e0{�e옚�<��Bu�c��J2����O�n"����ړ͏|�I�[�I�#C;�� �����听E[�����w+��v�V�2Q��g��%��V�?5���~��Vapz���x0b�=C
���*�Td���]��},WW��v[ܓg/��ˮפ��ddZCE(){��a� �[�	���R�5��"�IP��zlY�����j��1w�)�E��'�Q7��8�ܳ
	���l�,}��KR���\.��v�q40 {��):)F�/���������ѝ,�mk�sB�M��&ۈ�:ō���HL�b�I8i�w��/��
19��![kǮz��%E2��ٗ�Q��6d�Y)�_��_��J]ԈJQ^c�l"[<Kf3F���vN��=sh(���H�G�QZ�QO�Q��d� *U� �⶟L�`��x!��� ��&����
Ʀ�����E�p&w�O���4�&d��8ą
�6gvPP���ac�7�Uv�P�{|O��Ğ�r����fJ���ޫ��`}Fķ��h�����Р��g��x���¿+���N��}]���=)m�s^�ݓ�\ڐ��LQoֹ�g>�Q��Ҿ�����rn%�ȱ�R �T(ZԀ{"`J�p�E:Cu����X����mٺ�H���}9'��4��%k��zo�����[�+�o>���6B�I��2?m�qm%`q�{�6*\�w�K�*;lDH��nM,�o�9a��sv�����ϸ����|b�{��ax��U�!�v��Pp��xݧ���Q�1Y��-Ě�t5�|��ߞ*�#� m	򮅬�C-f���6�9A�Q�ZGuvPyWν}I��Ҋӳ�Q-,�l�2�Q������Ýέ�B�̐��Ӳ��3Dn+���A<�C�HM�ײxlc��1���H��=��ץi@�2��V��f�t2ѵ�ڣvq�@�~ʫ�an-�3Ō�P��?�4 N��쪦�]����>�!�����J�<�Kc��ڭm�)��Biy0@��+��/��C�IX���i�, 4s�n����%�&;/ǒ�/Q��?��wu�dB{Q�&�������sw����5sm#u��� DG������N[7� -�tO��Y���w{�<FТ���/ ��8��#N��|O	��;��K�
���ta�AA�+oġ;�d��:�r�UD�S�AS �C�
x���L܎��<7������z0�a��tUv�/(o�F^g��~Hw@]�ݷ�Ÿ����� ��t�35��]��B
���@#�=�t�6�/-�>����/����诖~WD�˭��&�e6a�Z8�_��Fwy�@��YU��&�Z>w��L�PN�:pN��h��Hij'&Jqj�uz7	3D�JZ�p�N:��ϊf>ij���=q�{÷��f��wS+��ئ�R���Ur�a27`N t��`��h�>���`8�� Q��)��0������>t�k=�L\�'�^E�1y��\S���l5��t8���龚��>��C���2T���{��#��ZV����|$���|�[Å�j3ˤ���4�0��L�g&���Sn&����Ŵ��J��Z��T�X�a(|l�sDs1R۾��=��vh��tb0�U��m��S(_9�a}�#,�ɡ��<�q�[�O�(�?`�� {�����Ս��+�����S�q$ҊqmÈ}�r�eB���W��q�b>x�ؐ��!	$���U��c؎C"��G�:8ОH92&��x�KsB�A�ap�r��ǆ7�+:t�wo5�з�لf� ��$�/�|�$xh���8? ��:� ��c
�*��r�.�p���<>�iJe��ѡ	6����f�r�Sr�sYZ'�H���\�&MY�����������$� ;۽�mt@�\fu �C�8ç��B(�r��o�5X��C��ZꡲY^k.�j���b�>3��4�X:�'������C	���*a���h��S���kd��z��3S)d��z�D��Jp�G��ZBe��:��;8����)��������cՍ�k���3#C*
@#I�6,���.?�g*�b�v9b��L�+�.��rܮ���Ҿ���Yh�
���� ��d��_��-�j�F��xӖ��}H���Q������Gv���v]�X���zCǧ�(}�rΏ�O1({��];7ga.�|D&ß���j�/��,,�W�Pr/AIs%7ջ��oȷ66'�m9C�Wo5�N.��	n�"��M����rƿ�%�~Y�w��6� �q���'�O��j�k힆� �ҶNߙ�y�f��/����z5�h{	5�lv6�����o�,}��yj���@dL�Z��3ʮ��o�G��\��r�Z-�Ӎ��O��Nl��+�C� {�F1�Ȗ�h��߁���	3!%��`\�]#(�h�&;�UǤ�����
b$�G]����/�QC	�͍����C��eb�l"�U��{L��p�E�@fAO�,C��E��N>!7�H%5���0�ˮ�3�dc�S��C���ǥv�\�w�i�3 jD�(|����ͭG�.�f<�|���#�q�	�X��y�?8������C��ͳ��$�OÏ#
�3������S��p����z	D�&,���2q����TR� J
VHx�!��qT�ݩ�0��E�)zKáG��,�N4��eL���.�*d�t�|�>	5c�	�@z��(
yAm�|L��m�E�@.NgN�覱(P򏲋��ٓ���75r��ŋk�=k<� ��Bv>vqP���\���2whQ�;�t�aՏ��@��c=�E���7;�<��M�q͂�^��=�A>BqT$4��G4�SS�;Qtckǜۨ�h��DUD���:���jZ�e�#����v�(�b� �1�H�Ô���,rOnj����y�7|�t_ÿ>��J�@�_E�{:�)GvA�ﵱ���|QS��!|"��
�9nx���Zp�Ս���z)���@�I���١ �e{�K�L��[RD^O����J��J����6U��vԟ9�����ԾB��BZ��X_u\����T�ԙO-;{VS��E�����2�^������'���[�r<���d�mz�5ֆ�4]�I*_�/j��A��%X�H*8��ճ��C���K�ǧ�E�u&٦�,��bR�Z���a9xM���
�(x�~�Ҽ�����������e���={
�Ӕ��p=!��V�v]9�tRh��=�~:.��Kݐ/�k��z-�!����ҒI���w�َ��ym��@�Kn��Q��.q�2��]�t ��V4�(��z��w�H�l��gJ��ٳ�xK������Y��y�i��M�x�n}c�D��Ȟ��~�F�=N��Ab��wA�S���G��:/D���i 1�)�� �:�� �$ϥ�߹1��I�똥��$:�����yܾ��h�f�����g�ȋ4@m^+�d�K&&1�3h�7Ӝ������r)�m�F��3��
��$(l�S] XT��Y�)�����������c���7p�Q-&��M���>Ё?���.tt�ʧ�s�Y��L:����	�]Z�\J��?D�
X^$�}�|��	b!sBk�&'t%D���3d¦����_c���?��F����1�ze4Y�V�h�5P�!ֈ� �x��]�{@p�P�<^�A�%O��OT�n�3���Ȓ�i
��V���aln	24=(����,�ß5+Y�@������n܌����۳cg�(��t�cX�e�(%�p�A��B'�tQ ��0�|�	TQ�{Ԏ�Ŷ�+ֿ�o?�q,hR`��[�!RLg�Ar-E�!���9���T���,���⪭�è~����_��U���n��-6t,��N*��[�5�(�,YQ� ����-����GA�xf|�K����4��,3�\io��P�śt$(�Zt@È`\��ix��8��A�z a�;g�F���z@�N�л� ���^ѷD
�%D�����9���!�{�s�N���!c<�[Ź? ��v$"f���!��V����x����`���-7���]��ܞr��2��Ic���9.
�Q]�K�%��@8WsZ����U^�F)���%, '	ߓ��� ��@-�X�����f*l���/Y%q�򠡮������8����/�`&��UV�#���#�<��~��Z��ϑ8�ݘ#!lo[��a�A+h���>�V#��I�ʵt�8�UҘ�C\��`�>)�H��ֿNsn9�#�E:��,#�/����"��E�Pl�z|���6��z+�vF�j �{�K�\ͬ��Q냵�{F�4Y�/���Q\�τ}^ׇ�a�>.�$:bb�S�+?�c�_����c��X�Ѩ a��w1}w&�\n�h����Q�DFL��s�������c���B��O�A���v1�BJw�K�K�LG(�������,}P�R�^>����y�QV�#Z����	�I��+PD���� �J4�3�4ȁ)ɩ`q@�m��Ӥ��:�f���;ړ�d-��C�պ�����s�ɓ_ۃ¶�z?U���}����`��!�D��)���/��!��Vj.��e���8��5j��s�d��;�Nb��&��F��lL4����c#09lz���@3g�8�Q����t�T��c�����!,9��^��=���&����y	������k���|�5ʙ�#"�y��������X>�E��&��-'��#X����󲍌R4�a�'��a,��<�v�4�UG�ojPν;���Zث���=b��V|�������`[�afZ]�М�x��+)���k�Ka1��������}�Q�(��4�k9tؾ��l�,���K�_H,��U�L>m��G�j���1{?������,�֝���{�eT��1ǃkO��j�*DNl�MU� i��5&78�GG�?)-/����Ĵ#�8MqWY�0�GKz+�P�)Oa���&��1`�*�p�XAĺ_��|8�6�(QQ��N<����_�#Kv>O�P%��j�;�q�b{|����C?+��w�o�y%c~(�"�3Hj����Ȥ���0�5f�F�p���&+%U��a!�pp�/�)@���S>5�+���nY{n)�eBy�'0�k�}�h��i�r�˼�i@gs��Ȭ���j�� O�^�I+%�$I	�V�u�E�/� ��u����X(��Ш`Bd������?XǪ���.^�b]B	�:�R�w_q��'�u�9�$�M/ȣ�d�~�h3�`.羻T&��ㅢh�Ȉ�t��u���`1t�%E�!-9��K�ƀ'�
��`���y�� ���ŘtUl��4�9���e � �V�,�K��<�_�@��@�B�=e��K�Q>�>=3��Īz��� Φ���W���Sf$D뒪�����@S���]���Ɍj�{g;�����*T�ܛ�'G�����<?�����5��}���k�n��Y-f(�� �G`Zi�ɘ�,�?:�f�̴[�fF���� 
	hCS��)W�ki�2�*>��&M�̦ćZ<$c����lN�Â�XN�PP_�B�����i.y�$�Y�EjX_CB�Ò�d�|�G^��e���h����x����A��2�Tc;��[��LVL�6*{���X
�4�,C`9x��>g�޹u�i !<
x{��#�1�:"���kC�\d�����6�.�ӕ�@��@C��:�$�F���k;��p���h%��Լ_�Zy������$�೼���=�1С^�	�N8.�ӪL,��B��Gx��)2��#����S�S���_N�f �]V�3U���aq����#���G�ޜ��i
��R!/�pX֩e��e�/����b���,�Ch�9@�V��q\ߡ?��1��Φ��a�ІH5O��`�l+�S���S��{�uY�0�B5n���n�}8QT'����&�2ڝØ`���/����E;�zA#*���#D���Q1j깤K��9׈�i����(a�zA]>�~3o<D��y���I�;�;Ҵ���D�m��6�BfVCH�ֱ���sJ�)|������
>ޜ�қoR�-�������A�觜�ù[�0K�Xٳ��ǣ����L�"��t�$���� ��6/zǸA��˖��p�=<�ރ%�DL#`n@YD��������[6��8H��}�A�+��}s�*��pG���/v_J�,��sw�	��k���%226Y}DM�a��U��s�H�B��Y3��� �H�D���ϑj��V�
9MEE@���Pɐ�MP�-�a}\^7cu)�I�qW�@R}ieK�͚���:7ľ�X�k��!�<���
S*i*C�t�Cǉ��d�'\�I���ive�����{���=�.�����S��*�P �9۬P�K�^��Ow��A�x�O��S½d-�]�����Q�T�{di����V�.R�9���T����v�K�>����a��z;F I6�5��nn)zyFھ�'t�L�f�U��į#��7�Gϳ[J;Y��BڡY����Ƈh��'��Ƞ��݀҃&}
ڼ�;nݲQw����8�x^{�+խJ�o�b*&l�?�l��o/��	
�Pv��@�U��7EV?Uo}�y��	2�:�v��܊E�GR��D�'�z>.��/��?��&�憉?��s�E�-�]�_3p����m��w	f���WYjַ��g�@��zj�V����
�(M�%���fՏ{��Z�Y��f,J8��8�r�\��]�_^�<0��$��p�<_�PtY|2���������G-;4���X�FFm!���~yp�`��8U �ӇU�t~��9�۹X��A����.)��̱���~��y��p��ig[��ou��,�H�mzv(�����w���mS#X��fu�VÍm�C���%�����"y�
X���%�6Mr��5�e��UY-m<f��}� ��2#�Q�v�0�deT��]��Z�X�/��dS�>�3^4 �#�_�>�W����u5�ɦ<Q1�M��ܧ_�aC�U��tC�e���R����w��w�'�o���S��k)�4�A�U�����Nϻb�����;���e-n��]�`��|k!�&x���M�_���Sp���)��@I���-��y���aD������.�&f}љ�����"G07�J�k���$�Z��/��	��`S�I��tf�L��uy"U�H��� F��|��z��5V2Gc�U.�뷙͉�>�_b��$	_!H3)o6�0��) ��m�l���% fϡz��0��)D���`����M~ t/M-��d�����Z���;Ɖ�ħ����u#4�9:9{L`�c�'��H�5؅2�j�]>�K��L)(z�}�W��y>W��mꅞ^���+���r^oC'Sd�
xO,�g	���A�:�7Ӫ-��)�I;��\�C�#�����U����$��:���z�kd��&��S�؈����0�97OM�.	q�g	Ч���Pg��[��=��]��J�V���{*�
P��C�\�f�]�� ㆻ��E���2�4�R�x�.x�0}`=9�#Ƀ@�gIl^s��d=i��X[E�\�[���1u8^���;հ�E2*r�{�1�%����<�'P��eI��#���#��s�bm�!��m[��9P�fKm����]�3��8��Y mV��"3	1���*Y�'�R�6)/��,��c���s�fz_l�4����8y��D�bG<j��klͥQS7�i�ۦ,/*e�PS\'�L��-�r��Ǐ�FD$���&x^Q���-?��\3�W��h��9v�t��HA���%T��p	]�Sƽ�s)�_nXO�,�%�E}D�KK��2��=Bvvg�i�������c�T�G8�<�ݮi�Z��B�9�9
�J.5�Q��hqњ㖦Y�R�}�J�!~������9�P������ ��:�<���k���=�-����l`є'�4O��(̧7����&��hYd�����J��j`k��d����L[T�;4.	W0 �W(���wGjH��w��ZM��c�����sC���>��V�p�BB��I�C�؊z����Gӈ$�%ކ�|���Kg2���G@+DԌ�F����������<Q�tC(4� �c�(F\TM�����5)��wT�T���r�!���4�G��qͮj�K���ʸ�G��?�˯����.x&��G��Y�����+54a>�	$�R �����"	�Nt�i=� U��W��~(W�5��/� Q:�(e�\�#������I�j���R��)��z�fE	���2��+g�p��W-�J�CWP7�	��������9�,K��:��BP2��*�*q��2X�<J��ҷ�y�]��\[�,��}(�a׈��p0�6�1�ao�8f,�Պy�`� #�55_���\���y�~ܞ��`CV��7��97;n/W�R@�]���ݦ�j�Wa:�>�~�?� 1�I�ڵ��'
��{4�㣌n�P�ɮ�'H�M,��6��N�Bh��Ҵ�?LZ�v�jm�̿�Ve���3yQ;,8�Db�c�bo��Aе��<B���v���?*�q����仼��l�f~5Zf�vO�t���L����j����3�{�qx[{���u�������1��=<	6�9��N��j�Aȿ�]�?'��ŻX��S~�{̳�pQ�YM�h���	���N\���hu�i	f��Ĵ�CB1o���ц�d9Lp^��Y眷U�̵���(ȮA��V�;�=E�3�	a�����A�c��r3x�ApLH;]��
�{q9�؟Y����G#���u�J1Cʥ�QT���5�B�UP(�&�k�	I��K��������[1Č�{>C�%�@��5oP��Š�PY����lM8Ȳ�N�Ȝ��ׄ�%��y�ar�2�f]�͹~%��|P/�q���
R�<��7��['�$./�K��tU��*��7����G|$5/��^�#�����H��Q^u��f�9�L���&��@Sq�� f�-V��@,�3����88�*���pɼ�dR���2��,�{���Աҡ[�GPŲ ��p}M���u���G�p�������1M=�&	���{��7�uWF3Y�+B��uj������ϲ�tZ*[:W���L�,�����'�1#9eK>��H3��<@�<n81��f���s�������I7�64��Н����!�ߕ#O#����V.��Q(�	���<�N�*���U��%+:���<o]'5��ߤz���LWdk���:��?ǽ��я ���r2[4K� Q}_�Z��2��Uo*��|���>O)��T�o�}�9���JsU�bw�D�����)����5
�ЅL7�p;��w)s�ȃ?�Vӛ�'B�R�����dOCs$�U37L�\���k�7��W*ϑ{�����%��{���ľ��0$��u+�E��	N�[�,.�O��N��_��y� ���;�l�Zo�+[nh|sB��aɗ�����w�yZ$����	��s}��@jp���xEuLd��P��Z�(��e��sTp����lK!��k��4�-7�9� �f��`�i�͓��U�K) R)��{#���D:��1)z���̋��r*o��/��h�i�ڛŁQ�Y������z�+�Ҷ1j�2" LU���أ�\�?;�1ZB_�`��⠦���*�
F��R*��sӊ�WZY�c+А�͝
���a�3�ʔ�$v_ ��-���=�wf��x���]�!;�B_x�H+��%��'AQC�9]+��zE\�F��`7�2o�Z�(������9ʾ�HM��-�I���i�§qj���Ua �^������{�;�������c�{>@���vY�<�d/&Whz)�g��������K� J�c��o��U)�~;'{�B%���mn�H��L�Ƨ��
�j4���EnE�%cԪk4w�| X6ʴ��-�E�����z�������r�ͭ�g��O�c�����B�i��T�75�����>tq���}ҎI�ܙp��-X��mز�-̗DGn��/r�����aR{�����o@_��5U���U�o��et�&����O�����bޞ�-^)t̶yK$>
����^��1ß$�Up����0���qZu�^s1�{��u�!��ܼ�A9�Rc�8E�xoI�P�� �x6+�I����^����
��rW}���J�b���p�	�ޮ���NG]��e���I��w�g��cD�6��-'i�-��y�[��U��p������Qlԇvj�'��l�)�ǚi�4�pa�O�)˽!GM��ʯUb� ݅
_�:J�.G6��Ja�Ig?r��#���F4�inZl����0X1~s&��A^��g�
c����	�@1Z�T��}���������;-����af��NkL/��Y+� v���eg�ƛ2�ߦK�b<��%1�j������j���I9Mwr����HJ	���y�m�S�Ә���s� ���?��z�G~��/nS*/Pɺ����Dj����z���C��u�S;�zC���3�K�̵���p�	'��7��c�����6r����b�+��j�����LlL=`T��1���8浓Qܼ�Rd@^P�3$a���B��ǖ��6�������-s��1ιJy���!� ���>go�w�c��`5G�lpz��APw����� z��S�K�U����=���BE!��4�ӷ�����M���9>����;����[�oy����N�glC�x�Cy`����	��{�~��V	U@�8]C���B���k�o�Oŝ�帨
����Ē��'G��7��&�+M�� < ʷl��U�
�iPY.Mf�Ly3o3$8�p�ǟ����tp�=߄Zv�qt�I�o,܌�YQ�f�t�7�CUg��n/݊�o-�W��:�Br��m���[�*��-.^�ວQ���4�F*�|����=|/�v#�E�@vg��9(Or!9���$�&���h^�mHT�[�(;4�-hƆ�P��t�3ٜ�����Low\Z�����~zs����$�,��s��Zz�RT� �i����R|��O�K	SPR�Ň��Ձ�C��эBL�p��(�Z]Q�mY�����؎�<��0u�����j�Ea5?io��W{�MF��CMm���;��TVu�I�z��i՜v@��l�@B"��Q';C��1b^����|�G��jSp�,�ény��p��(�N�[R�Q-D�R͌�h{jM�-�\T�9OB�6\-����-�1��i��l�_jHI�E�f]FSX���Lޛ����@k*o	�]�~���|N}|�X��PY����)n:;G��p�z�p��/�G��?$<>���vu���uQ[[*��ţ�?߮���T�&�
?9����}nO	��)�I��Ϙ�X�L������7W��_QdW��Η�m�����๪~x�D�b�4-Q��5�aht�=����DtK�F��b��}��cN?��n&�S��੽5i�ֿJ�&���(��Ex��ɩ��e��	%h�mo՗���m���ɨ�����(���lg�j[���g���5��޺�Z{$����Z�*X�l��b��(҂�� ƍj�y@#��'%|��g�I�����Q(3���;�
"�c�T!�#%B�u���d���_�;�<�]qӃkܧ"dD��r�,7K!��a�8�9�@�*f֋z��(1x��S7.u?3�t{�ή�����.��0o�>e�V ������ʈ���ȹe_�=��}("�`_ٌv�-<�05�

�a�;���_����Bcw���C�;gwn�4i��,_�o�rH��k��0�%*�^J��|}��E�����</r=jt��%f����!��ӯ!���zS�[G��!5��ڸ������r�-�қ�3-�ڃ���$l�,=����Ք+5� H	�E]�W����6�* FG��	����W�EB�6����o��ߝ��5�O�߲�.D�6�뉉H�DQ?C��k1��x.�~U�Vfk� ��Ň�O1;��D��?�W�����M�X�lG}=��ud\;N�f�	+�]N�;q<Z��+������jm������{sg�_p��F%Z��0h�m�ih�Ѐ�*��0��(�W��yk�j/q��(���q�('��~,b+�d�@B�vz{� @AC��9y�p�c~���W�K-ujq~���f�>f�2�Idw�Ņ�����w�u={8�3spwy���WX\��ӊ�D���7�m��F\C�J� y�� Ԉ��ݔTM5EB��E����٤`�r�?&������F���-5\�mo�oV�L���ë�&~���b�^�0]A�G}q]h���w������z�+{?nh"�(l�� �,!���wC���� L'�b��g]��� oY��؝u�n �ۏEo�o��(U����"�u�&�~�I�+�0wM��Ǡ��g2��	F���6=eR��kj��Z!;/�����q�'�)/�����HaK��߈[H��gp2�k�� �e��Ղ[Hs�Q$P�ޅ��t4U�8�<�
�U_-�rS�*�Ѽ���N��t"���Ip�
��t>�u��8:!S�EV�JH�Ã�礑��[%��b�����8�}���ɡ�e)%��8��۪�їO_|�c�;<����W����RL�v��S[���>�p��U[�@���7�^���{F��:#P.�K����i;��$���� ˻5�%ㅄ�Kն:�dCf{���`hJ�&����9a�����}��]���!�n��z�.���t��87���&ܞ�y6���d�8<���d�tDb j�JT�X�k���h�:�&�~u�eh�Qt�!1E��9�'�A������΅J9�r��#�m�E=XH�ލ����U}�y)w�N���,�ڟ�j��	��`�������I���\��<�>�7�T(�j˦d�fX6�u�ӥ:E�kv�= ��I_s��ۘ����+�"��k��,��#�`5�p'�JH�U��E ��
gi�oGt���b��,�b#�oE�z�s�Av:�NS��'F�+���փ�Z����l�lsi0�%��Aٗ�?"�ׁs�@)����b�D	�-E'L��ʤ'��h��p= Z�w�=����W_:���Tu����":���<??�\}/Kv�~OE���M�g�:;�$���w�x�h�[*�!��K��SP�V�or8p(���%?(F��J��;g8��ٙ��'�7�T�S� ��PO�*Q����F`b�F$F_�L���4�F�rNҲ	]��̹]��m��^#7/��/U���2|���A���l��|�x�+��Վ�5o`�e�w]��ZJ7O ��&g�CV�����W��R����^�լ�	������ȟ�e�~�y�4S�@{P��Ɣ�O u{.etgW2������K�^@����FC�a��T�$/���Ȏl˩�s����"�:�ݏ\Z��qVA�m�R���-;���y���37,SK�k���Lp�AXv9�U���4��L��Hz��X����r��X`�Ԁ\���mnБ�X5�Y���m�+6��8f����Z*@�#��̿,�X��	TK���2�zI>fLJW�X8��|�?����ȣX����dC䖎�^���(m[�{�#4�bD��,��T{��*��1�T~/�\��;bE������QE8^��9nk"OON�Y��qǒ��1ِ���g��xG92���d�
��X���*�����1I��H��I�����{� �ȁV�+T���gpӞƚ��2����N|�ţT�(��vq�3�[Mz7�����h�ߝ��N4�Op�*�=d�`d��mͣ��@{8 ��d���L�-��=�6w�	�����1!�^^����Љa�#�-�q����w��@?��8��'��)�O�@�����j]���'d�����ء��Y0+�!�.Zdo��R�Q���DW�L�~��h�T��x�R�M��)��KȹF��AlЬW����&��. x&��:�!|^삞�����B��`Mq�6BH�$!j�!���ɧ��r���9����݆���O�'I��P�EQ^��qa2�c����1���1oJ���5�}8�2�W�M9��0z��s��I������S"+훳E���a������Oc&�n���c���)����6���+if銱t��C+y��ڏ�	��ɺ#�#����������=��x�b��D�?�w������2�A$���0���l�f�sU��jd�����w[6>���#��M�U:���g�֚k�@u)a� 8P0��*��޻�h5_��-̀{�kt�a�#,�_�}�Bՙn<$B�/��RY��~�%ԫ���a�U��ۨ^97��g�RS� ���vq� �R���vB��젮��i;nwK��zW+�&	��d�d�2�駇���PD`����o}�D�V���~J2�, ����ύ�����&`s���T��UX���#;�ؐ�c�:N;x]rB��/��4���LSy���z����\�t4|��?�]g�����_���L�2q�D�p@Ղ �_�(I#���C�w���!1o���od�!O�G����ve�g�����$�WH$�y��'��y?:�ה#nv������}O鋮�q�vQ"�Oᦧ��C����T��+.>����N�����W�`�Yf$�;S��T��!��<��R`����4NJi{�ʊa���Y.�]������^MM��<��xuJ(�����v
�cm4��̀B'�m���k/��5:�2Rdp�A=v\���,Cz����-E?L�x�������5�		}�'u�\��LE��P�U�m�M�\ƿ�zԷ���#���uq����q�=��+Y��V|s)�����n�,W���Y�Zl|�=?]���j���vF���%KAG4��y5vGzs��\,q����R9�Ro�C�G��&������%E�y�'��0���ǣ�������J%yY�]�����7Ah
 ���Q���2	sx��U�.;)��Z��y4��H��l��E	�`f7�p�x��$�b�4���u�W�����@	�9q�Y���m�o����M��`��r��ȁ�K��2t�e�d�⤇Y�C�M6�.E�4���cc��&X��$v*nq������"=b�ϓ0{.:���!'��:��߇��Y`�%*�cgv�i�� fK���>�������O]6��I����|:KI!	�:�tڗ���-`%��ed|a"}a��Tu"r%=�*R�E�
뗦���S��q �,~wjy%�П�3A>u򘁨{�O���>S�z�a�6O��p���n�ۉ���N�a~]�k��nt^W����Uۼ��ݼK<�
SW��Ί�l�EWf#D���E(��Ȍ0e�Eq��ٱ�{�`6E�B��m�Z�qy�ih��M/i��u�i�l�?���nT���.~G:~>��(�b=��4�0���ދ�u��@pS!������,��7������{��.M��W����z}r�L̒��z�,��f�O��?���!�HJ4���].�pr�%�Tt �U6̣��ݛ��^�Hx��B��ݖ
$�Y��y�?s��;�|��k_K��Oi�{D����c��+����C/������KD3[���B�z�"��q�h��_F�۠
�������C�v�����Y��bߡp�"B�$ɜ�26��J�O|&�彫�߃v@9��_�릯K92k�*�~�1�Gq��Ғ�>�H�ja���>�#l��ؚk۾����tH��A�`Qv��)�lm6��b���a���k���q��'!��0��D�*�����Im\����.E�s�E��X[.���?�ؕ󞻴�lg7�K�Ӄ^�����̫�Ə�YA�'�~�,�z��E4})�D���^}M@�!�3w�f��0s4��ې:! �o���y������gZJ�H�9f+4E!�C�?��b h��7��}!�{4��_\!�{�@��z�i��ɧE*#��P�w,��n�3��E�AȑśJ�t��!�J6��I�F�'T������8v��Y��?�i]������?�掿c2�����Z�-�=,��zc=тV(��c�>ec�l���uQ20qр	�7}���(3���S��GY��^�lY��b��C ��#�	P�9]���P:.ENe:5��e��m����$�p���HWU�|�����|l'(3�!���{�Z��rm�M^G�T��]��Y��NM
%V&��/���������N�>��?յ`?�/W�P5,J��k`M<����Y���%�_�����L\rɏ�Z�#f�j0�bC�����$�(>�y��_h8�}Ȝ?�a�΋,Fqpt;��/�gYet>��o-�9�*��XZb��r��W��Ca@&�Õ�������"[r Ϙ�@Po��?�y!	���V��)�k{�LP�̗�K	�a��o)��+M�Ҡ�+x��v�x	��N�2O%}���N{��t)9�<�X��ӓ� �`��
�4�޺�ڡN�
�G��zj wN�D���L�3�t�͵cٺ}�Е�朲\�5��۽�����r ��G�~�)��զ��wh����9O��R��T�$g"��\*�%��H� 3��
5R=��+Xv��� ��-IJ�1�A�L��V�[��Ͽ��b��H'?��������֑J���;�]35�L6��C(z�����鷇B�4w�T�C�_�P��K��qUp����	��R@���4б�O�T�גvp%#5s��ZAJp��ͧ5���[ï���<sU,�j���(��)�qwǄ#�է����-a4f�8���Y�א����>	��8?��"%~��D�yv���� )i{<@�f��`�յ�v���zzRft8��r�&X�,�ג�Z^�����;��<N��Uj�D�v�e�@S�[`�MQ��8iҩk���������6�^0P�
$���awt��+���\�i5���@�W��N��N�ר��2T`6H �����~{�(��*�o����>�|���d���B0�U�qw�5��l��:��%��!�u6t{{�'��� ,�rޚ��v�J�
/�8ԣ�K4�6p����J���c��F��^��ѷ�̙g��#P,��8���?���'q�*��9�1*2!�]���ޓ��') N�JHX�Ω�tl.�b��{����P	�ܓ�tK)?��Ovm��+�b3ȤV���B��,�G-M��L\]��F.|�]}�ڱn�����o$�O%m~=4�A�*�>T�~� x�59;�r��T�*|��_�h�ʣ	���b�bַ�����W1%X�r��	�		�}���V�L����
�Q�����;��C��w�8�������*��z}���`�{Jڵ�x���@S0~�� �l%3��*�f��t���0���K^�M�+s�m�����@�^���+��,IG�r���u
Y�j����E�ܰ�Hp+�Fn���� ������f�}�����w��I�g�UCMn��,p���-�Р�?6� ��o���8�G��_����;�?|ay���� ����P� t�$f7�~��[��M7Ӆ�Z�9*`ꑴh���u�C]���Χ7kbow]�x��	w:K _P �	e%}^ �(UO#ש��qɩ�Cړ�Q��J�DP=�C?L��A6�H�5�J�C�4�R�6Fx�Hv�����Q(�W�C��9� .�>;����Jڭ�s�1R��t�k;Hs:|OB�I�M���z��x�)�N�hF$�.��p������8�J9Q(��*n���\H���I��đ�����xڐ9Z����F�O�{mPG��Ay�ى=߇.e2�������1�m�E�unq�����P]���S,<�W�*.vj�"���6G�L^���ζ���F��zBn��/Y�ˊ�N�'E�i������w�����Z�3���oZ���O"�6�ׁ�@�c�ۋ���=ej'x��~~�K;K���gj}%y�$�%��ٯZ^������=ްB��&�AF3��0�<(�d��9s}#Ʌ�H�kI6w<��VXa�_�)p��TK^�,�yh[V<��(�T6�ɂ\�RQ=S&�c�Ҹ�]�8�H�<Ѯ8Ysc#B�'�TH{����"��`�8p�Hj�]�T��f�<�]i�g0�n/���k������k��}Bp��ڱ�E(�΅@2����d��(���������h���wc`��lb��c��V9��Pz�"�I5� #��{��N�v�g�T�³]i;�Y�ˀ�Uaݧa�+g砪�-�l;���n6������c~L��oo�b��ov(��0Yo���S=�uv����P'�k���$>�s/��[
P5˟����F{�K��k �Wh4��o�.�}���)P��Lձ�ڥ4o/���0zD^��n.�xj4����U���g8`�뙺7+/,�,c�;+$�P�n�kC�TxaFMyo�_/������g���E����Ԑ}83S"j;�^FD@��SP�|�݈��u�B����k���`g�}Z˕3Y"�;@)Fy�'++��@�ew������0�9���?��b���GFK�/���9Ѱ�?4��"�=q#x,�R��*lX.q$-y
��Tf����P���QX�b��+�'�g�T,���\��g��+Kɸh�%���zc6�w��Y��"j��W]f�W���I	�b��m��D����i��L���t��
�Wtw�W���e�06����\��n%�j�������HR��a�K[8��,�T$�t=V��������q���K!��_b���3�m~���M�(�ʪ�Ԗ�4}BN�0�	���T9��x�g@���x:l p�o�����}��M~Tͣ��)���	~&.��z}����{z�D!p�}�E�������?I��G?�켏���j�|��u����X�n1�Z�quI�Q~�i^��s��b�	�$�X��E|+=&���y���bd�2z��(Q�#)��H�86�h�k1�|�3�e�gG6�R^rC�&���4�<�|�L� ƻZ��z�f�zƃN�����x-JK�)PR-Y����nɔ!�v%���g�	�/b��7�m�}�m)��ц<��MH*�i���}x����MM
�r�P�l��������@LPI����q�D�Nb�Y�����Z���uy��-�ט�@��7�����R�������̔a�ry�.�K���9RϪ��o#�{FRq�����C�wRu�o��,���(�巓�0�,�˔�g�W����q!Xh�<�N�6�+�w��'���CD����ٔQ��W��" 1Z��xʨj!�X����N����	nj#�p_������}؜^�#hۛ�k/��#���E�K��@h�w���=��pz�j�4��@�	��W@P�%7���{W�I��O�euU���GN�t�^t����qr�JlB�E��ݝd���p7�˾�]G
�ǩ��؃nʝD:Ҳu��,������R
���pChN!�;�����
�鰶nR/��^�=�W�??.�|�}t�CVs�sq~��n�(�P�B����"@͡�����۾V�b9�6�]j/rdt�(����_�#��3֖�1���p��#,H�rO���M�
�g�{X�+����9������l�.�pk�J�ƈ��d]���S�/���fB�������
~�v��-���}�ۯC+_h3ݽ��f�.f�'��*#��h��:�7Kب��_�u�͵�p��F�ԟ��?IKuԎ���JE�IeH�1 s\��(�����s����� ��*G��m	9�K.&8�PN��-dv`By��������2�r`��ݴ�Q��Y�M��?��݂ɳd�u��D�-Q�c癑tOH#�3N�hU�T���݃�`0�/�&�֣��R�"�����a̿ͻ {2��K
u!��p�EFf��{�	apj�i�iX�34[:��5>�T�;^����¯�k�V�E�u;�WG���Oy�g��x� >R�['�wI'^'+�H����
#�0���̯�-�F�=���W��/"S����y\i��عJ�EV�����(�$�L�'����0`yaX�ݮڕ���d?dn�%8a� *�μՠ�爔��U��վ��V��2����ê�pT�0�ϙ�XRODqZC�N�+��c5;���?�g���{�^�!���z/	ԁ�<վn���SIcB��m��GsziN1�J�]�ʄ}�)� V.���	ZC�s����ׇ<@��Bm�Np'y+Z�9u����[A�[|�@U�`���K��`�.$����&���=<�M�H����Oۆ�����������8A��Ǔ��Ϳ}�PY���?�4ĺf��82!5���g�J�9W�	1ɇ��^`����A	�ċCq}�}f<P�c ��_&6�>|�9}A����;+��9Q��{4|�Nv^Nr�v!ǃ/�����T�.W�ݴ��	A¿fS��L���irВߞ���8c�p��Է�6-?�'bN������TX���7Z|�^ch���GH.<�ǆl�(����J�h����1���e����%�k;J�]&S@�wz�
x�;~`Y�6I���Ԟ3牋;C���T&�(
g-oLπ���F�񨇦��Ȁzr�&�_~��&��*���]2�H�Pn���2bv/��ӣ��g�>��JӢ��@v����N5�����4�&��so�M���ǧg�9d�|Q2���
L��X��}��B��яd$	�o�[�2G>��R�9�����T;��R �"�5�)n�*�%h�$�]�����;�6�mI�W͸�!<c�G��M߲0��ۦ��Q˫b;�th�QL7H���kj���|/��,Y$������QwI�I@o�c�W;c�ȁ�;��QȀL��?ZM3%�����w��e�V"��C��h��t~lя���IڼG��`����P��c4��e�����U���%����B��R.�ݓg�f�T-nQzI��2
?�f���4�,��O��H%~w�QhD��zd��c�_�/ ��Aa�`y2�8�.���a�*SeĞD5� ð+)X#C
y�5�ۉ@���f!��"�7Gm�:�`������,��|;n!��b:�����#��~!D��0<�&����{Y�4�L0�,����A�s����2S��3�}����/{h&m&��-�.n���	��!�kH@5�Ȑ�B�H�rt7ÒZDE��	�P��A~�e��r0	�U�_v�AJ���5wGQ-��w�@�;���W��|S��}su��T_�� ��%l�x���v$<���r�_�	�W��Q�j�3�i.H��]~�d�f�YM:�3=Q����,��CF�1�U�Ր�s~>�����u��b��:���/n�_K�)���S�үr�}�t��g3U̕����ј�)Ћrȷ̚"YAd�������PL4u�f��f��4��)ԉE�-��uIL��E9���(F���Fƻ�ꫀZ�@��@��ai������AN��ǖ�W�(�}y,��i�ח�k�x�6=yP��;m��U
�(l��֣���ILc[�Yp�Z+q� �j�_Sd�Ue-O�6.��b��|e0���r�!-�0@��pͨ'jv+�x�%�8�K`v���d`2rp�y�A�:�ؤ���bH��l@���p�`���F�Ϗ�Lc���A)#6�G�0K{ؘ�!+���.�ː)fm!��Q2:��D1�����A�Ab�|v�"�Y�Ù�z��~;�Vf�+�g�:K��+Q�����C�%3_�5���g8ZF��q���M
���+3Ǆ�^$YQ�H����l��"�0?k^�ЋP4�e���`՚��G�a8t��KfL���������&V�gRހ��g����s̴#}�δ��4�K[��av�~3Ȓ�����Ey�ÐL�����L�r͇�'%{��Y��5��h{ɒY���@�`"%�	��|��q�S��N�q�Zo&�E�v�!�azeI�t:O=�w2�@
����g2�9�:(�Q�a�Ét����}Ҏ�ʗ�D �"f,**=>O�U�p� �ʠb��2b�)�M����"pq{ľk��.Ě*`\ڙӾe�*<�X��#����+��an�۳��,�ۂ�&Ǒ��ỜJ��@�i=�=�+2��%*R��#|�@�8{g��Ӗ�O�x⯋�и�ڥ�F����)��e�Z�0�-oqs�*�����Ǳ-,9@cho*�	�¦1`)Oy�߷�	�vIS���٣R),]M�͓�=R�)m�&b<�B�����pa���%�� ���7���|B���~���?�1X@ž�������r.��_�^8P�%�mg-��=��(��:�T\t�*(���N���z����%�?���2�Y��	T�������"�ft��i~r�<Mυ�~0F+Љ�9��.9at�2�>��RZ�� L��BJtӧ�}�z�*�T-~����6tM$[�.ic[�v�ڂ$[����h�Ę�������Fk�۵C����/]�AZ�NP���	�A���g\LBz��}��C�u5�����p�U�t��|��7l=7��8ѥ�j�B�P4�X���uU^�ΣA��bUw�֡��'��8���{4�����
�z�5�A˹:���*ˤ+nj�\V�=��H���,�RM"�״�l�����C�I���N��H6�b��MOTZ��W� w�G襢ky<�1�$:�ؽe	�t,*Df ��k��F9��@���3i�xJ 	$xy�
�`�B���D���g�K2ڱӓ�s�A�5$m���_O�xBq��泥~N���K����K�n`���wI|��vx-z�3���F�<	�9P4������������r�[ϥO1�6�*\j�3�.AR����)+6%ά���X��!�SH|\�J2�����=���d}�/�g�S5�T����ύ�d4D�(��֡�-9��Li�V$ؖv�D�T4z'�
�H�0�L�<�I�4��[?I�wJ���W���kT�+��PZ0��l°��5H��2�B�x{y)*��*(��;���e�?��@����p~&nl�{r��Y������b�Eͥ+�

�Z������;���	�<����wy> ����yj����쨑�+ʪ�?����S��@jo��4�g�`�|�h��7��� @G����k)M�����;�Jp�\T7F읭sW���{�];2U�� �aW*��F
�J\��:4����T5��"c�P�L�02'T���爄B��	b�P��������Ѿ�4��8{� h[�+�=*��1ɑ�S\M*�ƽqE�Z�H��Ț�ކg��Rl¶{�.WC��#����n�ՠx��\�v@��>�:���Q8�'�0�]���#(�3dg�N�R��߲v�C��9�6�8�OlV���#��A�*��h�Ep)�I*��8�%�m���e�O�Ĥ�6}: �a�u��d��j�>��ƩĨ�����7�ʄXag|�@c� !�h�X'״ݹn�����f\�e}�c)7��ww�w]a�U��R��Aw�,�~܂�{�T]$�y�Vd$bv�NQ���H����"EA{�Q�ť�u����τ ��hh#� �k�N�mS�~�經�%�y����]��N�1j|��u>�Y��Y�t|η���|�~wC���@k���g�Rn���D�`t?j|���/!��[�N�f�̝����$#�9���w�
�c�N��2�hxl�:/mW~�<랂O-�d:SԀ�+'k|_���?ա"��>,Q��,v �f�*S��2m3t�u �/ۙ���� ?�n��v��������ɞ���g���G7d��m���p��|%c7����LUi!-�Z��^�#�C�w�@���%"���H��Nρ�1��6����wf�Θ��=N��|��\��fOP�|Z���6|�0� ��w\��t}�����jW��Z���kV�J��@KY�㇟���\�B����2�e=M�C<�$��Cf�B�b�%r��f�<O���������T�-�Q�����rF.:�/�] ���X���Z��~{��{�LS�`R�>j���b�4��.�V�����ߍ��3'�=6����� P��f��[ꍻG�Np�iT��f	,+���S��6���~�E�%`17ol&ﱗq�R�J,_����-@ޮ�k��ic�������/�Jt�����~ ��G�[�����O��k���������{�`Ԛ�;��6&|-����A�<J��J��l3���7_�}��@�~Xޟ�/�RҏÞϠ`^�[D	y�̭^�%�h���z
������]�^M�tG�ϡCX���\�tQ@�ċR�wL>�6�\^�o���P�l?B�l�7A�!��>�X��fK��o��9/��~/�XW~ '��kF؊��g8V	��T�n_<��{�T�_��H`�G;�#<|!�����V󈥹ʔ�.��'��^���
���M��y6k˦e{�l�421����k�M����) :g@�5��Ļ��T
U���6�*�^.��O�?7��5�Y;��b2�E��w������y@�����z-+��Q)+p��";ѿ��Z�Bh���s=&ί�gg�?�%aAΐ��^v�>%�")҆��<X�K(���Oܬ%V~�j�}Enɸ}e$�n����G�)M%&BI�}�����<Q�t�o)Dљ�^�,�qbP*$33�P�˶A��WB2㼭�
���<}�``�v�Ezf��Nr���o0�.��=6��K�8��I�~H����[!0(�L��<l_]��&��o�G_������	��O�����P�e*ח	����E�D���7u��봕��}Y��i�*KG��Q��2Б���'�^{�Ot:�
����AYj�q�¹"b�8�d�"E54��T�(�����o�(��K� s��/ve��XF�yU���N�v�ғi����9��[����Ö9)��zaQ�&�ͦ�QߟI�����b�3�Fz��]�A';��ѱu��7�fH���f�@���^�,X��V9�lD� ��깼� (?�O����<=^fòvSύj���:eSq�2���)A|B��c>���t%|�sx7:��I���-/����O���'e#��3upbY�҇;t�w'L�y&Oܲ���٠�
��DA�)ʝjb��g������P�.&�lL_���?��~U��v��X�ג'�>��
E홸���M^�B�u'Lu��Jڑ"c���Q��f�h���L��xYq\NG��݌5?.P��I��.��(�.ه�ƿU%C�5���Z��(�BS�}
FW�/KFjJ64��o`�-�+�85��փ�P�j�|���Ӿ3���H���mu%Ղ�9wf����m0�(���$�llt4o�c@�]v�Py��OO��c�c��9�wR�a��Gr�	��F���ɺ������RV�%��x&�O]�����f�*�+����&��r��L	������b����cG=�_v7VG�|�͇G�'�3h܃ �=;�'��{k�<x¤���מPUS�:;�7~����R�F_�;93��i�|A�)�]��������ߩ?��������̢�=,h�i��>�n;��J/��"�ʲg�|�$����Aa�n���i���H�l��*�h����a��1�'�MV ��̓����1ܾM[����PD�"6�����ޕ=��A���HlA�DHD�z�}�ë�-��f��/�:Ra�X��>��ԬHޒ�������&0$�7[�^��2���|"��)s�i�봞!]� pi�~�N�	�:*�eg��A����1�x�}�}� }��J��-I"d�L��x�#�s6v�(�u���Z���v����Q�����9^�F\_LC�W������P��{Q���/,�gJW���d�x��x
�C���-y\Z�1P���e~���J���|Jt۝��U�%������I��񭣓��og�&�sx6CX
�7��{-y��
��_�F'"����k�n��q����BwU��jK� ��۾�<����WM_ �j0b���7�12���yi�Xq�P.�ѡ.ݛG]�(XDb�9J*3`��/�5H�_���h�
M�{Оr���������0��d�R`��m?�A�wu�Y�"P
DIͿ-�k3 �tB����5�6U[ d���0V�/)�h�w[���7�~�E7���a_����1��$��Z���\�����W!P�ЩQG8���B�Uf��Η��L��vih=��9��tQ3wSO�)�Jim]'��*.m
�Z5�@�ӝ��|^+'ǅ��Ҏ�����i^\%���`G9}���5�a*YR��UF��{�~Z�J��h��k�R2�������_j�|�#��K�`���cI���opzp��Vz*l�M�*�Av�ra̾� -�j��4u�[�2bKE�h#�����1��b[#=�\YhϪ���� .�{^��+�g�KEȋYTF������p�������W�h���d���[�Ki����N��8�����'Č�$8C!�J����1Y+�v�(�s����B�#^ ����T��!�s����=�a�cV	X];���k��[�φ�2���q��*�{�`��esQ�.��|��7�c��&K�<���&ԟs2�e��K|
㏄��>Gr�����A��KW��]ڄAL�T��p�ߨw2;K)�DK�slF����{l�V�Ω�G�(�B?��x��J��<{���� ���S�+�M��c*�䥀E�h��{4^�� �kMG.�Q`���x��X��E�`^u��؅1�2�V����֒���'`�(Uzh��W8�+���hu�"�m.T�2�N|1X����Q+�[֭2����4�t�V�)D8+2�q�t*�X�i/� K�Mw5o�ɚ��]{MҬ��A���㣧�0V	�~Q*4���������e3e�cZ�Q�~��6��7'�oC�w��4,���;����UH��]e��*'D�T33:����J}��\uh7?U�
0	�ݤي��h��9$����P��!��v�{Z�H��̌4��+���#�� ��l/�*I�N�u�WN�鵊�vƯ-1$����c��.�3[����A�~�9�:�l������PȒ��S� �ʼ�ϧ2L�+�{��R�ө����j���YJ-�&=?�L��=������Y"󰒸��b�a��;���ή�@�$%�^��S!�pqC����'o��K/�aQ����0���L����T��:�ZWʿ�khg*x7�k���0o#lQմ9��©����������iP)c)w;�n���e�M���DK"�r�]�\�8�y�𓸉ܪ�b��RJ[~#�Տ��;��7�--����E�91F]J�qa�(J�|�7�M� d|�p�_tw���܊^������4�`v���9�����z��4[������*�@�<�V��"=�Q.���(��B�x�ʼ]IXU��S�#ir����n�y��0����r7s��W�U�d��y2	�Z���.6��\�"����S�����)����� �6�����RCqW��xO�{�2�}rRXz�����.�`)�U���"^-�r�Lu%d��}ʚ����V>���$�L��y�d |,7˦X�� B��mi(�n���w�f��_BX���O���v��RNl�q �\但��Lj�`�Ҷ6���qY[�I�P�R��-N�Z�ƚ�|��?Q�w?�{��tr��>HK��)&J*{ސO`�E��muY�u�B���a����]RA��r`T�ϴ���70��c2 �1�l�
jn�;{fRP1a/JP�	�C��������n��W�͘<��/�B7F&�F������؂��f��R��h17*H܄��DJU�?�d�M�|�Ƥ���uP 7n��пH�+�����e[�
���>^9AIl��(��R�6_�w�����	����R-���Ѽ��݅7�zb�Mg�d���7��v?7���`�l�#�Vb?�s��S}��:z�`.����y<���֠����Hm�U)���K�mWvq.Ӽ������]��s���Z�⥎��ǐm���l� �j��`[��l�����
;d�%�b��ُ�?J�<�]�Qs�S����r��u�;��1�����:�\��j/M:E�����X�Y���y��pWн��.f���<��o�I��!Y5v�^Im��y��S� `�g��*T\{�E�@�B�N�9FDMIf�,���D�%�o�f���\4���$��/�[��b�nκ�N1�W���X�]E2GT�5����#���'>V=EǞkG����D�����7�Ͽ��!�^���j���6��V/�!�T>S�3������$�e���$��HQ������%t�jld��n����&#���!厍��kǝ#�Q���ge��T�p��V�\���Ă̜WOySK"�o�9̞d7��c?!3���j�>Q�_���v�����|�u��Ю�@�ŵp� )J��o|*˗<L2&I����J����9k�L��v���7�;/�#�?��?�?7��Q{H݋燂��3����Ãzs�^=��p�(t��yB�8����~��;|�?��ˆ�_=����fɁ����Y�c���0�\���% S��Ī��*[��d��3�'��EV$��B�������������\�N�����Szʏ��\`ļ����b[L��[�L���?��Joq��j����T��7�V �m>��"�b�R�`:5�>�u�}�
d���2`9�20ze���P6JY�.�#��J��V1p"�J�n���4������R�i��E2y[S��J�;��GhR��Uףř� <���|KIÅ�����B��f�x�<�x��.8(��'��-�.��\���,�հ���J�yY��7��bZrds�#m�U�FȀ::p�1IhO̣d�QY ޛ.��Zv��ޥ�����Ҳ�>\&�^����./�v��Zw]JjP	=F���L����<&�N�-s`��NA�������x�5��O���Z��5G�J��v+O�@�<��qU����z"(o�Tʞ���;d�Gr٠a^��{DA�����Z�r?�1`c�<X��c�o�n�ޣ�;ߨ����/v��E�^�r���ڰ(�c�����8����)�\��y}�v�7���eP�~HS*l(P��&CE�0�ײ��L��1���;;����=_���n\��qV��"��r�T�pS�S,���J�c<�\a;0�v�6��8ҍq��4��J�h�t����Ԧ�ɂh��4����������`+��ʹ�s��N�y;�zٙ�8���,v�ǃ�T|�	AŘ����봺@ţ}�K����O�"䬠&���,�O�ir�	{�γWVNg��vH����O�5�7�`���#��S#�~�W�]ֿ����Ѥg�p.����e�C3S�L��y���YO7t��+�}ݘ�l��D]��Q�ּ�v�Ӵ0e����t;���C��hQ��h�3�pAf��*�%�b�n!K��8fEP�K��D�ׇl������9��*.�G!ʴACP3�����û�zQ,�������y��e �2�T�F�{\��0n�6 �~��I��d+B���p^����t�'#N�K�1���ܩ���bx��a!�X U����<pY�u��Cې}�w��{]����7�H�w�i�� ��}x
��V�q��ل.,N�)y�Ͽ$��.��C�0��W��P(W<�6�V�K(��\FQ��\l�Kz�c<(Vba�Ě����nߝ���^%m&X�/�<[�=�~ �(%���.�[�(AKe{��D#>�s�V+]�V�+���Ű�/-��!�X6���9�2�%��9��<�Aqв�w��.�Kp=�rq��9��dt�"�1s��K���4{S�|��\5>�Q<��\����8������\�h��ݚ���#Y��I�WO]��1�ك��j
E�K�[�m�P��q��-Ӳ�윘��z�S�PN��m�l�E�_�":���X����ߠ,�OAl�r����'\�ԃW��c�ۚk�=�!��L�H}����m�)��f��g��dե,���&C�oP�k��2�Y�
څ��b׶d�	 څ�r�Ͷ����D�¦��#:PN��J{��H�|��'8����+�W"��6B�����w��J�U�����u(�b���#�zhw���������x@�����i�?s �,k��'�Y���5a=�g��s�5��B�v�h;{Dl�����?q'^c���[^������,=3�gk�����Im���Hk�v���;W��Ȩ��O�~|�&7�nԭ���ʝ�Sl@#����22�V��ʵQ�� �s �E0��u�նrpc����,��.�q���|�ޑ�B:�(.	n1|%�b��� ����ι�C���]� E0�C�)�ˌ�wɭ ����(�&�Cq��o}i}�C���g�E��!��--R���C�7t�=}��m[���Z��Ȩ��ch���� b��焴0���[�uP�cL�zO|~�����OG^G��_�D(�9mO��ioo� ��xE�>G�A2�֦)0����W��i˦a�z�3܂=5�UI�3���5��by�5�M������	�R���{�U�e����S	�q[���/�ݩ �ɛ�ra�t;4g2a��T�ʣ��Q����^��)�9lz��,�kgRM�W���1�3����]�J�X���=1��G�n�P�=����C1{�OH��a�����E�I�cՕ�!ԻV˷Q+�=ʦ��	�����x
6�ˇBб�<�gp��`*
珀#�{�i%d�fkY�Oxr���{��3����+m0*ڀ�=��D��w\�a�:g�����V�~���ZbT�!-�j�G�^k^���Ej�H�F_1��,Q���ls�@ӭ��	Q|)��TC���3��!	�m����/%��y�B����
�W��[�_���ÉujH�ԢQ�74v�� �~�q�쒤 B�2�����|��3/ᕷY���y>|��h��MH����FcY�f�!B�x��Ӆ	BՁK�����<o���x3*.j�L[�z3����[����	������Y�l��RR���Lr��:����3vl ��
53�ȏ��5��ۋ�����ᴳ'8w6��s �U��\�	l���� �0V��*���GG�ܐ�M#�/�P���̽D���N&���2��>b��Zf��bSR5��<jVo���aa�J�܂�L�8��]z@�Ǥk�!����� !�&��� ��V��QɵYb����-ďGb�9]��;�fފX�tŰdo5.Y�! ޝ���'<R�"�L�Yܦ@O�4W��X;�����KJ�z	/C,%2h|1gRfw�e&�s�'A$�&�;�1���MU��-��/�Mҙܟ>S�j3z>{�x�N�JgA�$�P�o��t_y������*"���ۃ�й���ZÄz�
��[��B�����_�����2ۄ��k�z���r��=�U�zB^�Ӵ+Ϩ�%��*Ǽo�qɕ��,�*�h��Ϧ�]�iM�#����Y@�@�-g@t[�"�%��O�@�lX�<ZQ6<�S늪���&��ͭm�fH%Cx���)�A��0���!򲣨�t(*�J��ˌ�$-?���*�ͧ$�n7-E��u�ӛ�"|m�H�~c���W��V`���׾w9L��\X��%���9�A]��-|��}5>��R�]4>����/Bq|���:4�J�SXzZ�VY�㮍��$���S�Tq�C�	P�)�M�TC�$m]���A���U��"b���׳�H�֬� zK6W1=��$?蓗�ur��gW�����سU��G~{��@�:]	^������XN>�"Z0��_�y�M�_M<�U2��G����i��b|Q<���ǑO����N�%,���Am����d���Y��#i�%s���?[���0�j]�3��&_��G���Nq��sa�܅�X�8�rζ1@|��Eu���`s4Z;}!����D�V�_*��{�^�V�5e)�'+����J��X�ʦ¥�-�Md`����
��8l

i�d[4��?�!��;����݅º��s3Բ��3��R�I��s���i.�5�;`���Иgi�ˆtP��N"�Ӥ��B�)�Q�x�E��f.8�����B�Ē���1��D���=O$�u��=��+��O3��_/�VS�;���`�������{#b#r-�B@���翑��Tݐ�5j�Q�Tv�3���[�L��P|���?أ��7�2�@s��I�������]2����)UZ�z�S�ށ�6�p�pݽX��]6��I��u��q��p�C[�e�m����Au�R��4�_s�j �( ��/�����щ0ڱ���$f%S$�
l��X_��N��y�D ��"$�}Ⓨ��Q,�� �2�aBZ���G�{���O�jl@���R?n��'W�)�fʝK�c�t+�G��lw�կ���ͷ2��s�qV��+�擎uo�ǖy5GpKR=kn]�^���,i$��K_._gϦ���)J�\����?(J_h����қ�{�=�XeW��+�A��ep�|��^���r��r��pծ?��7.�	��n;}2AQ9���J�  �G�z?w,RN�ݱ��U��q�<���w��̈zg��,:<H�i�i^:s�M&'[��o���n����9 �f<Ȫ��^�\ŻP7�u��Q$[6�����W�,$ch�s�D7�-t��M�#X��?�se�����D���e�{�j7g.���r	^�y|0��M�o'/�W=�EI���c�X�G��r�$0aUȹl$+�����:�@оT����.b��)>a9d��~���"1�k�/�s�AܽFQ۸9[}����ڥ/��( ^ƭ�����s��]8�=@)�E����~���/�l�����/ϜO[����F;i����Z�z�`_,ɑ��#�n��_
,�ב��g���8��2�� �N���#	nds��5?������K��0�V���?�pN�L��Q�
����++�S��6���_[�Ό�Rz���i!�m���t�"�,[����J��&��=4�#p/��b�:��\�'I��B��\�H�����R��fŭ6`��f��g"�ü�X�X��r���ӈ=�px5��s���,0���ZD��=n��t�j��>�ee����*�e0���`���T�x��mUQ����<��������Q>�.��������>U���m|��)Ⱥ&J3Mm��U����K�ΟJ�.��/f�!qf|:k������&�6z��sD��|�4�I[5��e��{��7�&�)��)&M�WR{A��eBS��>����ϵ��η!3
�^�8��q���7�nP�<��:IS�	�Y���lC"CLG�G�6��B�<�9H�g���־��-~'qa��x2t=��zVy�u�)�6Z��
R��m��L��W�o9��B�+.�4�YJ�'��@ҩ�u�YW��H��0мv�|ԅ�+e��F	)nM"&�~�Z|f�}s�n�]J�n��ٴ��_t/<�W�8;u�&��/X�8��F"�����u1�+��:1�����hn�;��fQ0�5�!�xP�-E2Z�;q��ll���踋o�	��L�<CŖ���F��\4�7U��aU{��҆j{�c�H;�h�؂å��)���ik_dG��:i2Ť+"ny^�6]8�^���\֋7�EO�u
r)���<����l��!�l��7���:>��e(>
.����S`�{RQ�Q<�C[ 1l���]��6��iu�@���c[z�.�=Vb�ބ����Kc����扚b��{�|�8'�	�Rt�(���F�Ay���Y�e����!�d����%�ڄ�x����ԧ��EI�~w@��6���-�ZƓP$�b���Րz��5!@�/�Ջ	!��XN�&�J�>>{Wi�J��nf���
��2���uLl��Ȉ��%h�d��_�Wx��f�i�ul�� 㺧:�΍3�ķ�k��Ff�����{!r�J�+�:�� *�Ι�P��C[�Ζ��|��˖��}̓oz�s�P�U��x�=����g� �������cv_�{��,����	�����	�ec��&	���^y�����)Gq��C����*-�����_pF�.�����a��[��Nh�`�F�p������*Fօһ�N�����8r��@��Ufqv�=[ĚBAv�Z��%6������Z��^&�Vi�.�`�<{%UC�̲�N�M82��)�O\]��P"�і�BE�2�o�9��FȮF�p[.�ض��ɋ]�a�1Ђ�dQ4G]A,�7��ϰ����XԜ�
I�<�"}���N�_[�?��b)�%̪gݔ�x|S>�2��
�z#*4f�5Q~V��5ȘO �^�^��5-k�g-�_3'�B}gСe��V��/Vj����S�[`Jpɢ6N;_�P^���LQ -'�d6��=m]7�z!Ww��КR�-E9�K�üc*PV!��A |�%��I]�1>�q���"~5~������ؙT]��tA&
�;ɨl����R0�������d��l�H�AM�����JM+��A�W����KT�d@[U^��	:<�^�kUӄ�;���f���"ʞ{J�÷/c�,�(-"+H։�@hE&��w�Vh�i��y�5����>|�e��%6R����ظЕ��VD��i���` ���p���_���۾#�3�籲�<�z7.�ީ��PH3�I��ѵJ���GЊ~�r����6��ǁ���s��c6	�T�s���Ax��3:��&\,��H�1C��j�F��[�:�3��-4��Sh��N=�r��^��p	
�oHC�j�h`�Ǘ� N�A�j7m�����\���w���O����B��'t����Ǫ?!����L�;
w:��V�"����V���f�Qf��>04P~����s�.���/�/�e���iCR��iX��ow�2)s�k���9)ш��G��CF"<�Pnt|	����!�s(���hf������**G}�n��g�B&��i����=6|���v�F9���(t��+�q��#�F} d-�c���Z��^�=,{�9���Y^k�)�{�����T����̴H�F?�i��"
߭��HX@'��Q�Z0���y�b�I��ՃT]B�D=
Ć՞�4�d^��"��P�R��/R�Z4z���ې�M�����(ϋQE�GXW����<!E�$M]7��u���_�;�Ih^�p�kR�y��c���&�f��º��1SF1��|���5P�|��0sZ���R�c����ص�ј��e������6iJ�A��kh�uF�o��I�[fF�7�׀%�8����KۗyƜ}J�[iI$�Xg��	��啽��M�ͤEm��lb?���������@3�����rCt#|"R]���g.����q�F�|�a���\_^�Fk8����v�_�L�h���=��k[�?��n#i�Lo���Q*E�q=g;�M6�vﾋ��s�G�vJH5O����6��mAj�¬�a���.:������Dr
]��:��/���bN~�B�\�*�z\�Hc5��7$�u7�R��h�%N�1F��� ��J� �q4[5��;�X8���K� ��3u��&9s�yG��r�����T��?0�j^P7���g�v�NH!�H�<
g��l>��,>�O��MTZ�`EK)�A�6xȶ]⓪��̚�ׄ�>h`�k�;�z�X���fI3�w���w*i�i
�/�ӐH���S}�3D�x�U\��� ɭ����ڳ������RM�:Q�F��LEߔ�:b;݅��iihݹ��:�~(ф�̀f4�5��V�e�e��]�l��fl��u��0���5Y�hQfj��R��`^�za��0��H��q�-����C˗v?m�l��9�M���V�A۬/D�S<�T�Y8A��f2;��n�c�E�z����s��!��~)���R%���}�A���)P�<h��g�`�ĲO'���"l�3Ӣz\	V����w�ε�o�����p�ל��J8�[��a�[������o<�`��n9W�k\HJ0�[/��F�,ؙ�/��a� mcpԵB����م	��Ӛ�� �����~7��E��V~�'l��ԑ���|	���(�UM�ϛgn-���
��v��#�i*�쳣����*ZQ��|�}��r<z�����Ѵ��r��V�F��xx�$���<�C) o�Ԗ��4��Ά��1.������vQ���bb��V}^ǸY���a�� `̦m���2�v���c��X�F
J��s6�J�\�=<S4ˁ��'W ��"���:�Y[]}�vS�֔c�Xٴ)�e�$�E��ۍ�W��fJ���Bo`�����J�+��
%=j$y��m-&���~o�����;
"� �W}�Qgrf(v�����r�g�ze��*Nْ��k�~�3�Lk�>�T� ��5��,��j��4`���?B�2�\'0��5!�"��A8�z$@iَ�����\7:�3\��� ���&j�'Mf神�kLR]K@S����|���	���g�tC|���aH�c�`,Ց�r߲��5P�_d	�9�7 �"�1�oOj����mٺ�י��A� Oe�|Q�c���������c�t&s�bo��j̘���]F&IQ�nm�Fw�D�(��/�1��b�_&�vF�nK��Qq����1�1}l�"�p�	�1q
�����C�'TU&G������Iߺt���@���u��mV�������0�b �{�����,��g���FN�Q`�?ĵe��p��\��YA�}'�U�@�f�ɜ��1b3d��,;�{f����x� �\m7�����C"�](�=�����!�i9�IO�,�=��ҝy��ъ�M�����Uy�>��6w׬�J�k� @���3W�=�-)��aH�{v�Dس�$�l��_��]�S���IJ�}*���>W��`��`�B���z��_�!@��0����\���MRb�LJ�Q�����ϙ]�S�e�teP�>6w`6 ����kA�(�`��&�+	��%�}�w�/�N����k���wg�v��Q���̝��+����Ϩ�qv��g�/��_�P7�گ���4��4˖݋����<xr�6�k�ԑ���޶*���������]{ML"S<���/p�,�H�*��M�G_��x�B&H�E�Wނb��r 0&�x����G|-���r�67����tZ�g-U��T�c	�tv���ߛ�LOo��$�ņ�r��^�ܛ!Y���d�3ܛ9l�<�^�{3�� �H���o��+����V�Ɗ�� |ڇ� �q�<����'���j�>�E���ÕY�3T|��]�7�����F'�Z	�;(�_��Zt� ������&F"k5��W/E���l��d��b.>�2vՎ@6yt8g� ���2kڎ��ד��3����q��ծ���l4j�3��5U��Bm4�g����]�� p�d�C��NI7��rUw<f�L0�_1oL���hM.w�k}��Ё	����YR9c��7��{AdA�_xS��f5S ��s����Xt�04�p `[q�n�A]����J��\�61r�4��n&?|�3)xD�¦�3��\���Aӳ�b;��Q��
:��z�A&�Kҡ[K�"��a�m���*=��Mn��%�'��?�m��ø^w�Rg�IMBL�v۰�p��\"B��9�Mw ��k��ԙ��������J\	�?��zO#6�.�{fDf>x��s�z���YF~X7{cO�X��%H2���Bd�͑A���w��=�Ք҆�R9oX̙��g²��ʷ<���wϢ��	�N��vub:y]�I��z�F:eθ�6
�㯛�?Η%K����`3(��O�cµ��a�==a��!�A���K�s��Z�6yth4�).AXV��'
�	�\������'��W���B�� 	����s�W��R�&����($��BE�¿�Im�L�d �^�C��|�7��Xڽ���[���`e�U�*䃙Ƚɘ
�8[�sHpN��b�t� ��&% ��e{�Dg_�F�� %*.%7��
!A�=�p"S筩�.k[�_8^QnZ,�S�F�Hd*�;��Pk�>-��ݮ��1�(-�	��D&��2?}@��[C-��=���&�z㓧��l��eѹ3Ȓ��R�a�Cek�Ԅ����zk�J��5�Oj��hJ��]U�k����|��>*b��>\���6H8�Aqg�d�oQ��h�c�_�����1]��-�C�g�O;
��KF�A&:��2T@U�I����32 �B���t|��;3�4���d7}����a�z��/G��#�}��Ə@-���(�i
$$#��z��L8��:��@�=�sS���=z��ı睟Y$�(n�&��h���zk�ͰZ���߁�u�ނ�p�;H֘��^nfAIpˢ(���Ԗ���=�l�p-��ZF&�7Bq�� ����i��r��I�y	z޻��"K�}Տ����B9�5�;k����GJ.�y�����B��8ʨWR}#��#���N4�Y�.���o7�R՗��P�qk�~��FS�'��/������5զ�F�������F*$��ʠ}��w@L=T܈C$��`�����lFqf{�J�pw�� G5�>�����Za���[�����"'I��E���q��:���BӪ�h���+�^�[�-HKMθ}����'���b�{�Q�`j� ]s�d/��G:!6�t@l����*Qr�VV<?Q� ����C�n�@wy�iI�Lî�_�Z�[��j���Ww�ocw5� �v',��Aq��kꫯV�t�!onC�tq�c#�Ogr�S}�\��j�,eP-]��eJ�ч	/d�y�4���K�0u'�>�%�)y
� ���3ni.]�Z4
����X?��=���ݢJ��E�L��DhS6w�4����,8��p�d<\�D������G�6�F$��0=$@5Eȱ�^a8�[�\�3*�)K`\h��p���ęh�=;�#��q+}�FL�'�,�%��.e"��Mg������\(�#m�J?����s}�YL�eny]�(+�`�fD܉��)3c[kk@_�'W�"1�h��ht����)~�V�u��؝���qT)��g=oy���tG�0����TZ�v��>֩��,�1ʠHl��|�����6�Ė�IT;|M��X�]bPK^����+E�~'蒈Gؔ	�['�8�K��(�<�^X�SD1	G|�w��aY°~��u�`E�`eD�������@ǚ�N�z�4/�43󑇮kKuM�X�o:j�l_�Cs���Gg=��V�)�����J�S�~��߱j$oKD�Wވ��ޙ�H������zj?B��|.����
�
 �-�˹`sR���s����a��}/IQ-
���v���aC_�>��B_���2�)Ѐ�:yS����24�l��9�YV)�1���d�3}d�5�� CV^��̒��t?�b�@�Κ�zE�!j�eU��\W`�@h��z�K'X�UoW.�p������)�jj^.���!��v�<�u��d.�,3U���Y����ͬc7n�|��5��\��I�$���f��#f���B�NU-�:Dcw�&NA�`�oN�;A��̈�ޣۆ�*��v�P�
�2�F�jQ���<���@�����YX���<mE_��F��� �KPY����o޹��-<x=e|��;W�j[�"G^X���5Ŵ! m'gl>���=�\�{4��X�cSy ��H���6Y��^' ��@AE���0;�O�L2x�?]K���l���n�I*�jz�����]J�m�^0���Pa�MS l�d�c��J�&�C*y~���Y���/���f���g��$n,�L��25_���3玁��q_os٥��:�e\m���o)��%���c�Z���RЍ)�N�Zc�K��E�g� 9�7{�ە�w�q�������Hڂ�b5�_Ξak�)d�}����
T`@�:��� �%�	�}���z9Ȩy�
����7�~��!]'���NA��{�0�HȒ�/�
q+E�3mK�3JV����� (T��#�[�PI�C���m�MV�&	�-��n�%ZH�,Fo�4�L��k/b���5�L���	QKN۩�ц3J�)����*�0�� �ڵ;��w�@��e���T���{�	�ʮ%2Roe�
�'/N6�Q�2R�IS�ڡ4��'��^�Ɇ�ҁ��pFFǒ�pb �l�W�t�:Ԯ ��56(X:��+�.0x�B��Էp4l�4�� �0%��dsl�̽�^��������̋x^��"�Y-��0��1�!�q����*K���[��&+��ŦT��_5��Ch>8����X��cbz��*�X��_%
CG,W�1?�iN�;��Ks�
)&w	�<�b'!#�B��s���KE0T�q9��D��*[�K�p��&�l�`�	��1d����<�����<��=�=�*I�p���vm2�'rO�n�q���6&t������:���ԕ�8Ew6 b3��t�o~�~G	��C��{܆`��Wu
GQּ~"�m��z]h���?|;�3%JI�K��-i�eIS�T7�g���t�3H�$��E�2�/�P_�Ȫ�[�_�&��Kf�E�r�/o�s�f���X��c��Q��o�O��$��bG6ك��n�e.u�XS���Y�EW�"?����`,F�}��/�DnL{��7��4�(J7���Pʀ���@ƅ�$��n=e������m��7#a����ql_C�(";q��f�������̂����7�a�<Gs�F�;��?���v��B�N�^�H����)[3�ng�vu��:�q�~�O{����\-�f 
�M:�O�ܑf�M` �A�[o�c|>�������)uG��/�e93�G���+8 y��9��6-���r�?�p�����/�(D3~�@ۙ+�n�RKUy����������\kw���)#��*�^
�����E��"�E��sAZ�*�rj����u�K�z�iJ_v��?�D�s�v���ܳ���2�~����!7�o���; ���k�w�͜�|�@�����)�mR�`F�"`zt
='��Â?E�q�L��CGL�,YE�>;��cθ��޳�����vQ*�
��OS]�N?�E�6��oy��b!��� �S+O�O�fA�lN�>�ch���kc>��'�Km�&}'��!b ؤ�X��J7�0��nh��$\
7���`)�D'�_�����w��[�cƾܧ��侓��k�XQ|�H����~��ש�4Q�c��"̢e�7�\_hu�C�Ğ��+T:��c�^������F��D�Hݭ@i0�Zj�M��W,҈�0cx�_����6�A����;nڽ�\��O�/�b�G�J1��ۨ��e��)��G�#�3#5��K$�<:X[ �F>o�w�\J4�I��3慽 1���ӻ!�ߜ�:9Q�u80̽�-�k/k�Iq_�)�K�a">�3�F�:�r7�v#@�7F ���ޭ�|��%W��rv<�Jє�Q307�g�����x'm�����k̇m4"k!9��o�˟���J(�,)�[{J��\yT�d������@s��H���@�W�o������E�+�2E�5Z-��࿟�2�Ó����Q���v3�l���\��1(�Wd]��P�B��VO��U7�w��,qKX^XDy���D���Qz��thC7U, ;�P��r��y�Gs$�9/ -OBLu� �S�����i,���݋j�?#�e�٥��PZI�1����z6D��cN�tQ���T���NCLH��B�iY�^J�-��[���"�>�j��g��pr0M�3�p���5Qv���S�������׷MM�,S�+�����N5|k�wݞT�F�A� K6�O��&��TpL��'{o!�@���ߐoW`�Ɠ޳�&KFX����,�\��|s\M{����u��yP��U�$M8����0)5�l��,g~�p㫩�d��{t��"1��q���]�z�u�v�V+���/ݢ�$�u���oL' ����޻����R����"�}+�4^;	B��!�����<��IR3j��吡+�>
�4����9xU�����Y�Ǧ����D�Ȧ�W&k3ք�s��m���'�7}�2��#�>~P�IY�"�#L@jT&�4��0$s��1)��Q1��8��8��렖���� ͭn9K���Q��m���/�����c��d�3O��*˄~�"ޱ��b���մK�y\Ʒ�?��A�5��[5]ҝ�PY�ў~�TǪ��1���z� ��0�?]�PTI��)'b�s���"�7����K��x~J�������3H�p��O9�Ĳ쿾Ņ���"��TZ9\�����#�{G�J�S�����F�܉��y���\�Ӆ7�(J��މt�����ҠD�)H4Nhh%sd�y�l�J�Xo�⎊���.��wz��W�cJ��W,/��Įԉ�/�mX��m`1H��	�B\�J-���Zɷ��	tR�P�o0nЙ����&���[w��핹�\4����|P��ͳ��3�y�6���ڗ)�(�p���ߵ�a~J�2���>��'�_������l�6��풵z.]�is$���p�B�ք�Óy-�.��]���J�87�m:=s�,I����� !i����|���-�<��c���V��ϣv�`E�ez�0�z�����,O;�0�<_w���_� �$�#O�7��Y���3�$���S��l���@q@�{J��A��p����5z� �\+���ۑ4�>P%L:��:|�*"6I�8�P#����p�6m��.4.�</+��(UT�A�F2�(�v��q��޸�3�j�."�ı�8��&	�>��δ�V(TI�������u(譓;�x���m�[�q?�(@Ҭ\0���S�V/m!o|{����gu���c���Y�h:�H2�����KЪD�E��Y�1Α��Y<u�X�7O���[��l�n�����P��E��S����qm�Q� ��
T�O���^w�֫�fsFlh�H���G��i����}dZ",K�<|�T�u�{*6M�â*�!��-VR�+�����C�ѱ�C�R�o +%>�]�x��� B���g��k����^��L��Dc�瓁cJ*��֭�i�K�!UM{Oϩu��P�g�ԑ����wjk�n	3gB<޻M�i��Pb��P]M\���SEa��,aγ
*��p̡I>`^H0�@JTSm;������Ȧ0�;v��v
�+ݓ�1�8r��l�W�N����7i@��Q��%|�My���&��u�_#�ɹ;�'}K��9"t"|�¥c�-cw&6д{K9�iE���s%_sU [����Wp�v
HH0p((kZ�����Ǎ'�t(�D��w\�"��Cم %�Nw���>|mw���k������)�Í��P��h�R-F�gc���)�Th����x./���i��6�F(4�9���?�LP�v�t��t~"�� P�9��JD?3d+��/�V�������Fm�tC��e��>��((bv�L������P�.b"r�]/y[������乘O��荫��׺�.���	kcM�^��`*�cm�p�dZҊ顋.:[ʃ�k��6�hax�R���u�s�k�)�<x����^��vq�j�Wf	�p1���J5��J|��<����:�Hw���%���ކ��L�=����9������:���掣��n=��nviX���l�瞒z�"��2���AoF#ӌ��_��sG���!y�8��>��Jݥ��w��*��,��x�A�G���52�O��b���Ȉ�D�<�D��'�d0)a�<����>̄f�s��@�:b}[�93W�:sE[��t�0H�G58uU����H1�����A2f�+�>�'b���jk�ߋ`�$RD<~�e^ϊ��\�5i�A�Ȉ9����"��� 2��-Om���ϋzgAzCk��Q��ҁ�rt�c��J�q ���0�=.:�n䊭��Ҟ��`��u�Z�I"�s#��i�%�L���w�X�+�I*�����lߚ�i.��ۏ�Z��KĂ]��<Y�[���V�`wm��h����ɲ`DI��{�B�v��o+�]�ʵ-��6z	i�_�κ���P���c3��[~��V�Q\�=q2����j����|��6Q���&Y�آ{�+�*��W�ס�A�Ѣ�eg۞V<��%�����[���!@~�s��B(�?t��is�5s���c?4�u����)ی6��A�}�r��8�A��xM���
e��O:��'0�	.�'��=�?��{��bl�"�ܻ�0ѫ�+!���:`>�F�b�y�����#h�Ǵ�B>���̀����m��� 4�|�M��u�X^�/���j=�m�(�q~׭eC��1^(������� 2/�	��kޖ]�	�j���Q�G��n�߅[��@���2�W����u5���\������~K@� �޸�h2�2�(�M�V�W�g���2�j�kM~f_����V�d�4�G_�V�Q�k�aamM����V�����[�M�fP�����t �/�X8�Yc9���@0�WgNW!�	[��4Ը�@���MI�)�KM��3� ���l��?׾�(��xG���o;��2�u�-s5�f,QX��J�����x��9n�r���������Ø@"��1����	u�4� �лo����Q^�w���/����L�����8��}>��&�qݫ
N�,�;�7/Z����w
w<��v=o�f���p.�����VG��J��iY��G-Ѷ篃(q��M:sX�N,���ʖ`X�=Bsf�2ʖ~��Mg蘻��#�b���߂���N��2o5���爡_�-���@COiT�[ NY�"��d��3���[,'��Q���b-���tK%2�0�W�r�|%��R�V�R��rq��ƀ��0i�z��^B�<H�2vk�5��c��	w�@��B|��o�X��>�����-���NsTg ���}�4%�t�7��1MQ�ډ���p�D� W:�A7{Xꝗ$Qz�䇰�F��F	7/�&��U���6|��ܚ!�+������<�ޞS҂X��k@6��� H//Sa�ex�8:�-%�՗J�}��6����Z�)f�[�8��Yt�3V7�ԑM���f��9����4�rt6����y���㰉��	��o ������G�AX��V������S���pPj딀�I40L�f1�-f0V���tT�Ɖ�k�����d�e���M��xR"���xb�v)����>�1�3�ș��KK�6�b�ˉ�	�$�M'�Ŝ�����i����Vx1���L˿�Y��'7��B1l�L9W~�p��g�ޯD�U U�E��Ogo�Tʸ�6�^'Sm�%� ��'���70l4+U�<����(��];�9��&�^(�;�#���A�����d��AMd`S�[ash"�9�;�3���tY���� 9����:C����g�xJ�<�Z�
�E<�*gu�&���$F���La�[�瑅K�����&��jZ9R�_���Ql�`���,Xl30u�TGoYh&��aa�2��O�G�i�7s"�
&� �+-�Cd8��+胵��5\��)�=���>(�����`��|渖}�;�p\���2�����ڴ`�h��0�Qo����������&/noz#��$�C8sɝ<�����Ꮡt�<c. ��c:�����C@�,�\�­F�ݮ�k��E)���|xZ
G�G��=?�������o�L	��}��G���b`3�:N
u�s��٬�8�O�,6BU���X/��h��*���C0ČOr�w�}i���=#W(��ܕ����d�VQs\]Wgϋ�-Xα�KCKf���L�<G
|�q�[�R��ϒ��6���Heڻ״��zU>K�4W8�U}��)��J��#$�����4 ��nD<�d�|�����YI�F6ե��O~}�vZ>"E�	n�(s�Ii�u�K����F�z|B�bSRp���'0�.�7��\x���R ��2��"$���3u')p�D�8"�6�Ai]	&*ixK !��:��t��T+�D����M�J�ѐ��S������q񷁊E�0����P>�a�+�5 .d�o�!��7$h����y�N���C�r���)ԩ/��1�>
6�`6�(�&6{H�36��?,'�;ȬA�tхqמ�J�(�N�A�� ̀�,_51������9���;�|� 	j�-/t�Y�$_濒@1\�(�Ń��2���:X֪�rϖW�Vp���e�'_�	��L��������	���f�2'܀g㲿 ���l�%������=4RF�`7
�	��ț��_��]k��,�c��l]:�=G�ۜ�=��Ƭ��&�S�5���&γ-�;
���j���.H���wXoCBVzV�=^�k�������#$RE���!#T���j���W�.Ѐ�~��Zf��Ũ��-j�d�:Z�E��#Ľ�W���1y���)Z����^\���]��g��л`|��S�����&r0@�V�bp����]����HR��K�ʱ{�IRklL��2��|+�C8�q�$�m-��M������ժ�|���w˶O�O��� �a���O�u�)�E�#��[8�օu�
x�^���SK)��ŕ��ѐ~Xf���H)�K��{~*�ݻ i��)w1��]`c�7���j?g@x�&M['�0_)��x�ǹH�%��S�5�o������X����/��8[�A��`��)�Tl��r�V�'Al��XL���603�C�k��]��ʑ7�D���;
�������փ�O�� �t�}��U�	]~�0K�\�ǹOa
e6�jF�tS��?k���	�rd
�*�"�����Y��}s�\\p�	o=7�v��k��S4Y3O,h�۴	0I�mˎ�K��_3�l�S�qe�|�v#��[-nǃ�@�Vp()�Z���r���7���.b�}��O����I'�g(���a�n��8��v]�rHR���.-�+�����Ǖv�\��!_K�:��s[R��&���_ٻ�3�����4I��,U��n#9�̼nc�B�e�y���q�7�����Wؒ�gn��<P@�Dţ��n�:F��r&��m{�k�uޫ�3�<:�lT|e	@�g�G��������FE�
�D�Xrge���:.�?Qnq�tT�u���'��^�ZFL\�!��L<D��@�K��g�n$Ez@{۬�qު\�Fg5�����C�Q��F���=�3Z��z�L��P"l���Ϲ�K�8�J��ڂ�m�y��+.p�3Y�\�B��to��/�YR�t�>S�O!d�C�͡��k>��$f�
	�sv��Ʃ঩`�CtƩ�.S��~�s(�`�l#�%"�?9@�MiXǑ�j�:�TlJ#W\ �]Gn�d�#t�26]�T�!Y��������L����ϫF���{f-x�.��+Y�T<�� q��yY*'�q0s©'�9��` �2�O�o(�+bH�h�K����� �������"�U��d�:l���O$�luaJ�}갖��`��:�kA��c ��Bi#zDᵆW v���|�)(�5cI�P��y���j��k��Yr���� `g����=]Χ}"{|�\���Di�<��K緋�jW�E��"�/���ؽ
lK%4��P
��Y�� -�lW&����\��!��(@}����$9C�Y��c|����]��l���6Â�v��l>Օ]ݎ�A��Q/+��}�eT�&:�#��x����u[��>״O4�
D��*m��ْ���W�:yYg�U	ֽd�x�қ����+�L�Ko� 6^t,$?T��g��=�����<�=�� �M�ًbH7����	��z-��W��<���"o����}ȟ��l������*�����뛙X�º�KL��mm�|��qD�ʀY����7����{�M��`ӿ��b56<|�*���p>��򁪰�2�˲8�� f��}��a8�k�4Ԗ,�u�pٷ},̋��W���
�G�O�~���OkE-7����(��Lh�sE����t3z���Bs��rV�hl@âEF�|�A��*��Y�4!pdo�wVIL�\�5��{#v5#�!�co�-����6`�n��ê�Kq�y�1�͹w�26���j�&�g
�C�<�l6M+P�������i�=#V�!�z�
G�至!a�4���7m�O�	LR�ֆN���Qa"H��V����Y���t?�|�.y1Gyk�_���L��nLcZ�e8�Ftf���J]��0�m9Wb��oD?�q���Pdv��5�e'�ǂ�!���z�������\�Z[�H
�o���QX���W\�6��	�4��PA�B/}�xI����_�J&�c�kly����ϕ���^=s�l����\��Ӹv��y�j�"?�N�/<z����RGc���T�ym���6tgj䤕�t�u>&q�F��hp!1�狤�v�ھ��ڟG��D�s^��_�7�_���2\���+���8v��R<�jݿ�g��h ��]X�p��f{��o��Ne��ǔ��IQ���BOk}�n��0�q/�ǩ���x?���l�>��p�������B� /�p
��Ѝg�2r'uPU��&�]��w��Vʑ·���bp��ԘY
�RV~�o��߄��Gz�F����аc�x���{�]�����I���aO2�(�E�鱛���P6Q6���=$��O��s�o���o���z}x�����b� �t�b4�W���J�\���n}�K�'�p��զ�J0㬭������dyV�w�vd[H?�o�75�}�K\<RmS�p�<	�.�W��k�(�c�
����j�M����l��5j�Yl3�9w�C�*rܲ�b�zm\��}M�Nz�D�'4�O��=�U}2[Cg�����5
�F8�}��*5g�\a�l��:���3�ڂ�iA��÷�[�D޿	����Č�0S��F@�p���lʀkO�ۜ���1��+�� W�y վ{Oj�އEꕑ��,�wi̬ֲU�hF�k�Z�!2�s�n�����$c�͵d�n�{3�W2�aPK`����<tC{�]x�w> ���n���!�֜1��P-��K�$��b�*^�}��l�	Q�2��;�A&����1m� *�*�QS��02�n�������]aH��ͽ��~��K� �{>S����*�;�%����D$w���C�Kq��GL���i	�&��S���sb����8g�UX�#	�F�א{��=�_��bZed:鿦�ְ%){9���
{%��_�1�}Fr釱���%僆�am�YTJ�{8��֞&�sTj[mF�����>�am�_S��/�gX4X�Y[O�]AvA��-���P�k���܊��:��uԿN�a�"����$�#	 ����6�m��Zi��4a74�6�-YR��ي����rE��7���S�r��yE�S_���C�� 	o�m|��3�5H5��[��ʱ�0s$�H9R�DG&�=�Jy��9�e�(Rp�Ӝ���C��Dב����o����{�Q$��
�#.Գ�C��;�N���h
�~���ǵ7�d�`l۹��߁7�_�卧���mxa�.#���!J���{������WM�;��30M��6�T��9��G�,�^d:���M���5Pk��Ʃ�ߗ-=�8���ɄFMN�ft6���?�Xĥ;��&�Z{F�B@���Q��X�����>�	[fVФC�[;or��[���7b���2�ނs}��5�1
�jM�=��`l	Z����V�
��x?j{��j�o0���:���v�Q�rM`9Oɨ�����[<tiYHu^S����:1?��k�Gy{N�J`���`��t/�7Y�NY�հ8B�#C�ࡩS3��xp�PaM�����i����c�|[#-_x�X����rN�AS�P�z����{�6Em�2�aV��6��s�;�:0u+c���f���;��;5O��zv2�TO�q�w`lEN� �|��Y�c���	D|��(�%(с6�e�ꊪ�&��h=h
+���0�3�(�{���N�D�ֻ�zt_���a�C�ʣ��������n	м�;�]p.Ȓ��T �V�ټ?ǹ}τ���W�,�+���K����M(�a��
�0f�V\����|8����4u}5�+���L?נA��y9���Ɓ�H�|YhV"P���?M��)��5c,i!<X����1�g��I�"[���7t9�'t��
l_�޷{����(#m���(_ǐ��p������L�3���uPA�����E���5KL\��[V��#�u�cd��;�Ҷ+;�Y65P&��;fơ�UN�����������vs�r��(�)Mi]��6���t���y��2���ȉwg���B�i�J)��y��{�<0]?��DXh#��n���x��1]{��~)�c�v�rC2|�".PΚwAJ*mY�L�&��Ee����u�\F�~�~��u����yqu��w�8�  �!l����]�H�z�{�R����$��u�`P�k���4.�v/�- v4H^����c5DUV%X�k#!�^���0���Y�~�e1gW:a�}!�'Ss��\ĦF@ZR�пR�����/��n�����Pkk;��#+��Ռ^Ӽԉۺ��#���f�ߚ{VD2QD�a�r���:�_��B��D��ٖ{.5Y��zh�1�牚5�K/�s���,���FU���:��#4�C��K��A^�Nl,L@c�	�%y˻R�L��J!��\���1ew���3S.ɵ���.z:�%���s�M�Y�r�ͥ��i"v;�\X��k�#ܻ��&t�UT�a���og��"�z�P��1Ԅ>�����9ܕ%��"�A�+厫G:tZ+��
��K	{*늊*1%8Fl������rf')b��=5�Y��M�Cs�h��jg/�c.x岰�_qqzi�=hG���r��҂�}Zz��-թ+�	+���,C����՟�zp~G4��?<�6�ZK��)���!(#z'w��y��Y���Ö\�v~���^������TN^�j7��9�5Ȅ�BW�Ţ�zLbQl�#���G�m���@0J��
�)�R��`~�Ԇ=g��9�R��x���C$��)�kh�d���T1@���tZ��)�%��V}'��3'�S}^�S����D�jb�=1��i�	��g�Wt��`k��$��\�kTt�?`h�Ǖp'��+������i�@���u+��.=��j��k��2���$ξ�*eS��inu��_(t�xY����ma����S��<�)�4�-�f��YD~��2W̎|�澫�ϙyd���f([]��KV���G,ZB�F��\�Z����侥�"��k_�X���M�H�mf�g:�89T����2@�3���R������5��R���<i0]f�X0z:p��`��l>��.����Q�>Jl�*���sΨ�_%�W.�3CPoZ�+S�����֑^P�Ʉu��fJ���0Y�P�ۢ��ȿy�u�P�K��+�G4��G�PC�j�V��l=KX�mOB�WaO9�(wF�$ү%�TE�4�.����Ә��������I�����!L�����%��>�J�� ���iwd; 鄽��^���2ȟ�CQ�@Ņc�[fU��s�nB���o,x��#����� R��	�Z��8�_X{JZ:�^���L�$�5�%�/��JQpk�����1�wKe��������[�2�$��k[�h3��3�i6ӊWK5;K$:ۓ�i���lU�Ka!�.�l����� %o�A�w�kz]ϻJ��Mx�'"�z:Po���U�PB�kg���	�?j��P���*Y��X����`39��.>ry�T�Ԡf�?��$�wM�=��+X�[N� �͢�GY�	�i�J��+
���4-�4�Y�(��k�<�����#'R���Mf����i���9����L���΃(7�R�}"0�U���lUX4�]t�\% �Y����˿��B����F�����]5�w!�ʳ<����U^(d彰hA)��ٽ��H�0r0|�ϫ�me���/P���`rp	j�P`��nLѣ��\ѳ@wSJl�����pb�&:���!�X���W��w��
��+����qx��3�݋٥�)�7�2|�p�z՚.�x��(*�(7f��!��|(b��8���n��Q%���jU<��S7�51����R	��t�pJl�=}?�n������V��9�,�Z^������ј5��r5��,ؾ{�P���)aX �JM��~3O�X�����bl5��C�Wmg6�4Ԗ�5JLO���IۖV3�-�*,?�]K��~��m�\���F�|�v_�`�8µ��=���		h��M�����h�w8�m:x��:%�8M[l&�a؄�;5ﺺ �L����9���^hQf�Ȱink�OWf�Ԉ~��
�Ԉx�?�@2�v5g�`Ysݿ�I�ix�M6�q���_t.�4���%�kV�|@S�'�=&��J��(�����0E��z��U��a �ɞ�<�&daA��\:�{�Vp<���ht�8��*��0��R����<�EI N}L���*�K�yͳ�D�\�����]~d��x����f Y:(��P�Ck\�썮�g�p�� I�j�~db�n���e�ݾ�C��J�'I�O��z�������͹����_��,ʑ��V�;��)����'z���$��3�:�� ��O�9�� ����9l'?FP�K
@��Z:���:c��D��m��Y�����$OCS~5}.��c�ҹ�
t{]�U�I�Ҡ2\}#�j�?g�ၰ���#!�:�o�S��1؋����ާZj���F�����f����Ä4���z�[3ŤW�^�ޝu�?���/�c�������3��Ƌ>&X�7�$m���"qM�_��B�h!f�NO��x2�vC��5���珙�SX�Q��E�*�qڋ��SChy��}ymS�5��g��Vv� t��Ū��#b�F����8㿫�6��8(���Y�4rkE�Uj:��<�)}�}l3@h�X$��(��7:���h���p��x��)dxc��y��	�.���3�\��c�i�y��S|1ԭ_���1�Iҩ��V��=�I���N���fLQN{��.FyHk�K��\�Fŭ%7�'?�nWI�3�~�n�7(�_'��H����l}�E���������f,G��c� ��܇���l7���V�n�2�7�o���h��Fւ�ߕ���9<xz��o�-F;��f�f��|8M��wtk���(VB�i�P�8j�ٍ�}GG��C�8Ƞ�(Ksmk�2k�C��g��v�ŋ��b@l?&S�<��u��C={	����N�[1p�S���k��"-ݻ��/ػ+��Pfp���e�ј���KL#��mp=��S�����N������kRr��$�6e�g�� /��s��^Ph`x�<��D��9��y��e������t6+�� ^��*��
?z�~c�7c��1��S��>�p@�ݍ�s��L&�����m��Y���i���R�`��S�Z�6�H�𘹆�������;cKr���u�c8@�\��^�O�5���Zج/,��1��ߙ�⮘��I?���Џm���$Uѩ�aC�ڗa:���4TǃH�]È�Vօt�\w>��Șjxb�'�\�~q��4@��+�X�"�,c�k�5���j5/�L��K���xQ��i�x>�a7�$�-.�X���Uh�zf����R*I~��ـ�}��!4��� S&��9b��X^��4 `���C�2~u�����F�*�q�_{�I�t�n��à��;��湗���#3�� ���z��*N��2u��U�^}�Z�~"t������1�>Zgݘ�Zz����̜B�8�_s��	+�m�A���'���:1LU|V�5�iY����&��`qH�1�D�lu���<�؛O�QdVw���G�!��ؼ�c�+p8D�6��^4����n�b<�A�?�Z��T��'�@;�?o��T����A��x`����-n���X���=r��`��粵��k�*y;qG �h��R���	,�	Jm��,�ݙ��?V��.��>�7ѳvŶ���G�%Tf�J�w�����v��?�.~F�
37�ڮXĄr�bl��:�	=���4`67��|
�F ���m8��e����VL�)�u�� A�vOK�翊^���«�t�A��]VR���.��-f,z��u���i0:a��s������6���>��ϐse{^Ն#;<2�H:{�9�x,����Ҡz�	f]�y��f��g��k�E�l��w
rV�)�D�b|T<п���q�\S��hK�XOEAK��6w>��IKHI���t�It��!�3�Ñ��2��Eأ�Ue��F^�5<	+��JC<6��5|6�8|���.4���^ڄG�c��n��b�k�Ym�������Dt�l9c�S�׋)jU����P����#�~��Q�l���pWk�#D��6nzī���$�w$�a���.r?�w�?^��� �yKc@��A@G�J+|��.������Z��J�t�< �%��Y<���i�a�҈m��vt��*�[�-|������O^�'H�j��:���������w�+)��z���/-�������k�Lh�6@��xb�j'���n�B#}���K�'������Ȏ[����za(�-<#Dw� �M���-_;����	�{���V�
�����[:��W�V��i�J�ə��<�W�=_씹�D��;���� -L<��!u?s��}�deWr��|J���F����(�:f���f��*�R��,o���x�^�H�|��ʔ�?�F�(�_�0��t%t+�@�)��u�������� �D�:�S` :J���&���M9%��jFM�xht�^Zᬘy{��C2�����~���F��d��M��3gf�J}�\,+.Ҝ��B��+�:%�C"������j ����Mem���iw���J����0�k 	��;�-���Lk��d�ߟgu��9�x��*�������Ym�#;T���?JL�r�?��l�Gf��D�� ٱ�P\�H�4��D�)���  y�%]4͏}����f�f�>��H;E�0a��4����#訴�5��a��W�M����7W��0ت�T�,����}�pHÐwA���7:2Dp�b����uޒ�8���j�+���N��i�-��Ň��Pt���^����G���Kf6"���Z�h��QN�gNI���1e4G��4�l69����=S����+!7�*�����v�嶁n)R�3�?�>��C�ɦh
t�ͬ��-_����/����h=��[��#��ݘW1�� �@���6?A*=�����~5����J��'|�x�s�Qw��"e�����2�i�l��3[��(�ς4?��ʵ=��NY!.ǆ^��*��b$�t���[q�KJ�}�Q��k�LX��.f��T>S�4%��s�?�_�u�-G�"b)x�V����gD����ܟ�=j��{��AT�R ��qbw)�h}
>���ѐa�)��=�L ��4�c�"8[$5;H��%gЇӎ�������>	%�}�sm{�n������n8��R���p����ϸd�CK�|����.�'M����h���#�Ptjrb�������d3�n�Y���:<L9��<��+��р����/����������EY!"�|�V�YM	�k�.7nG��T�<�q�x#g�R,yPIȲ��Cm&V_�_<f����j9�"��Ą�A�-������E�qt��L�2��u:L��ѫ����]�����ș�yV�u����3
�T���L�P+X�-=���2?qw\Z��G�=GF��8�j		�Th�0�@bt@�)�HR1Z��i�_����5nd�Gm�w��RH�*r���`i ?����q;(�K`�U���a���)�����#� ��~IE�v�1D}F��G��P�+��ʥV�XJ����8r��f�T�V5ݸwVr���4�22���|���l%��v��ti�@@�������@)��*ڕ���:T���S%�n?��9�tƐ���ȼ�_	�,�l�7�D����-Ct��qq�Ȃ-��ڡd����^��
r�o?ģG��R�K6�嫇�q�r�[�9K]{g���ufΥ�m4�ݾ�0��4S���� ��<2�~� ��J;�R��#�g�xF"��*}(�>ڰ�Q篷�稍����$i��D�m��l��.P�����YK��5���N!#?��I�S"�U�<�Ӡ��bB��5��K\��'���n-;�=�ǔ�����r���w��W��Oxy���ps�o���>D�Y�0�?G1��p8
I ��w(�T\Tݺ�}��ܞ�Bz�M)�i�b�Ȋ���L�pw̹�ME�Xʬ�T�e2	t��;��c�^���u����{�B�ԙF���(��=H�)�K��љ2t��^N����yk!�� ��B"�>�ci�s~u���☐��Le_�rP��k�/������@՞s������+����e�?�zhr��<K���xa;���p����v��5^��^9⻩[P� �����亵`_����^��S�x�b_�6a�d^�S �H�\�=X�v����~A��3�xk�1���_���FkݷL�%rw��!��n�*�,����&����E�E覚س�p"�I8ЅC�7h#�-�J��J�V�T�ΥUO�J���,6���^HpeJ��+*��Iä2�I0��Lo�b6�g�u�\��ŕ�ip�JeO��0��o���w�N-u����a��LT�.���p��6h}N��_�Cz둥X;��f�{9hƕV��:�Y;/%��U�H�K!��I��1�Fs�k��T4)k��.�'�X%��%�����_dgW ��0Pʉ���s������y�Nӎ�e�\��'r�;�[`$�=�C�1��r�8[��\ 8#����bG9��߈:)# V�����V�V�-Q7?WD#���z����0���ohTO/����p�j�)!tIT���=\�\O����@��%e��õP����z�,�ۼI�Dn��[�#$; ��2����?��):]*"f��|�kv�qܓ��T񭷏_��j��a�FQ}�__7�;j�w���t�@����.
��ۭ�ز4�ɝ���W!ynL|��zľ���=����̚�����u P����ʽ�߳�+��56�,�׭��"���!5���S#�d�?j+���&�!����=:�?\�:a�'���#O7+�93r|��ʌ��j(YJ���;�O�|uR��ޏ��J��i+�jO�}���u��'��^����h�zEK��Uh^Kr��M�j�q���+�����t��������l%Pp��޸��Щv�jT�6���/�YXY��ڧ?!�	�� �d���X�� <)��9@R#'𡉓7�^�t;C��e���0�|��#�d��t-�l��3"��Z���v?��`�¹&e>l�� � ���Z¹^�JD�f6E�k�-8΀(É���ǆ7�.�p^^(v[���8�١�N�
UⱧ��x� ���@�(����
����{`Q�23@���yqG,3P@�~�����"m��՚M�r�.�o�@G0bގ�y)Nj�0
?�x1�]��b�0�����Z�����ۃp�#^7 4��xkn|-u�Q��ս
����wGKL�T6WЀ}��7D�9�R#��,�Y���~e7�;A�w����:����Dx3�k!9������ؐ��j�{-���4g0Ț�aq�)Xk1�����}�V�.�%<�MRK�Z~"�-������dW<��S�89�]��:=nG�iA,v�y��&.���g: �I���8����yK�����l'���9�Li94n@��!��"�[T�s�D���.dSC��c����U�}G�;�9�{��,�W���������@7V���REv?(<�(y�*<ŹFQ~^B�^�R � �x7�d*S&�A��=o�I��\�0�+��k�a�3٫��s��Xc��q��$���H��������f����3�s�E���S�sͽ��(�w��Хxx��������BBZ�O�DX���<�w����b��g��~��W�bEW��a�X\7ݿ.v��^�؀3��W�̐� kyg|'bvl�	W9ګD[*`~rChoY����|���[\{�n �}5��X�n4��ϭ4�3%���%���֏l;7�����-����Y���'�-�@��#js�Wѳ<�W����M����̐�����V^�� l^��˂��U���\�3g܏�F�O�{�TY��)z�|M����I)�����$^�U�(>m�d���������6\�`;א���`������fCJ�(zsAo�9���$`��o�B��6��M�k�j=<�le��	r|K�.Z�Mq3���&�
����x�IM$2�G��E�]a���>>�����?I�&d)j�j0���ۛIT�!'��v��B�Q�;�N�iW�J^��p4�(����~�VR�g�;�%�S�PL3���"���]�մN�z�Vܤ�d�$j�w�$��@��TW����9�e�	�R��s\(�6�rסڠ�X`U 1�F ���NqySlCwt�o*�|>HT��ħ��Cd+�	�c��O;,�@q�%� ��w5T�����6j�#�u-&�~[� ��!2Q�R�? �~#��BC�d�po��VO���w�TWJi�}�k&LP��{S���a�pݥ�y���֮h�"QA���epC���;�:�q�,���%Gk��p��Џ��5���! �ЬH�Y���0�¢����{U�~s��-��zo4����Ę�x^p��b��>�Z\������}����������{�<�yfQĪX7�/{5�x�D?7�A�?����i�~�t�Ν|��4�<R9)!�X�l�%
9�B	�)%'��U���wlvP4�z]Kɍ��$�s����_����mlb���#Kc"��;��*��d7{P�)�QRl����/��ς*����FZ�D�t�Q�B��p2E���tRr���Y��
yQ!,�#��+����&3�*�U^�Y���^����J!c�h2�ޞnhv�������$���6xS^��.����Y��Ի�)szCH���^Mx���._�w��(�ܰ�����^�_*�-Z;�*�,��yD���o���8���)�l�[�;-6������iǏa6��<5�TB��'m�Fc\����J�.��"�`EN��)h77ɺ�Ǩ�爉��ӦI	���e��ܦ��N��������N�h����e�c݆�����K�F���ŴQmF��Ǿrd̰`��C�MߖE#*l{ѻ�ŨA�ƶ����l"5|� zXJ�Ƿ�r�)�y5D��G���G����@PB@���|�t�J�<0��.H��YfU��i��E&cҗ�6$x�@�W��h�mu�E)��=q���ʹ/�{r��\qCQ8�Ae�,����V�[u��7?�YRm�٘Z:�q��$U{	(�sϢ9��K��'�s ������i�^`�j5��cJ�����I��'u^�����e����C�g�˿}@-�����s�*����g�=�~�_A��D~ �d���N+�0��((k�U��&�^������dvȄ�[�=��I3e87�n���Ko��~�����C{	��8��Q��I�]l�p��k����6]�~��U�]���3�VX���BV
t����xn�TN�����lx���!�q�o*C|��.�sh�ѭ��b�^������厄	~)�9�k�7�0����Qk�o)�#� ,��[��
׸��5�բ��}�ˬ tR�{��g�tr��u�'=y�.ǒ���ȉ[(A̢Y>�:kCD��a�w�9��c`��/�pRy��W3"%�W�~��9�W�QԈ_�����*9�4��9�BUȻU��'a1����Ƭ��9�7ʲP8�7-�H�ϰm�뚂�)�6�xM��/���#�A��|C����ۨ
a�+ʃJe�u�d�ʶz���
}Ŕ�îɟ��bk�b�W�����sM���u�Vӆ��)�y�v�����u/dg4J��0�MI��f�_56�3Qf1A�T��ݺ$�:Z�w�OsN	:�%"]i e� U�L��T]G�F�b�\Tb[a��.���ͦO#��q��N\�E3Y��	I���8ߎ�sT��~\��2|	?�'���rN�@�H�e3g^H �����K����������WJݧC3zӽ*<s3��$?��wg��c�=API*qX��9�	��wg�H@ys��U5g%q	(}G�>�n_������+��(�"���#��slv���ƎDT�y X������䌤����+d�˩���Gz\M8RO*�G/���sώ�C��^�r�u��6W֧�Ąx�����:����<��,��� ��J�)#z0�/�����/ �t�v)�V���%�u^Ⱥ6N�8n�F�:�EhE�؛�`aЊ|uGw%ݤ������� ���M~�9q#{����_@�n jANb��=˻���Q��[ZDB���'ľ0�����+	`tde�Z`a�h���o�g��	D�',ңb��fo7r
�l��TB�ES�y�{�M�(�!��ĠPH�a.��[�x.Ѿ؄��Aׂ�ٰ����,�m�ެw�`IFTO�!eo�E�_�����V�����G��f��.1"�;�3�
X�(z�b辄����,�����8?:��k�ua���Ǹ[�K	�pW<y��-	����)���p�Wg ~?N\������I��ZXZ�liML:�d6A�[��i����t��������mhvI��,��K�Nv�;-�m��y��c/�U��<�L�O���G�&A�\���V�8�ԅ�U���-n7�b�j��b�(�z��%<L�29u�ջ�v����NF=o��L���2�� ���lYņ���v�>���o���8qW�8^U���#̟�-WRvA���{1�㚸�y�g��u���'(i��ߺ��dϦ��<lz��l��ň5#�?u �e�j��ց���F�5+�^��|����-�m����8t|ď�Ŭ?ށ1�ʊ��@���B�̔Bmo&���@tQ!�0�*J�t�H����Az��xՈ��/BޑbҢ9!,gR[���߄ ��8�
�q�#@N��&(���׎��	9�x��p`ż�q�����i~�GP�V�ě���6)P��닔%Un�.��J�����Ka7�f�D��9��oc����?� S��h��]{ϰ���g;D���a�@�OzlPh�rW{��2Ԍ_���3
�^'�5���ȶI��
�Au����}�`D����K��kKOP�I�o�+�۟���lT`�?8A��l���}
$.��R��5����īM�7�F:��>�\`����o)�oI`2��}��hv��NtU6��5�����*

�m��~�V*\ݓ����}_�"���&��O'm?nW{˥�|�g"��i��'Iܷ���H��ЏJ�(q5�,���{	OB��m��K���*yۉe������F�W�:����$,�f9�{�������h�
 �o > �	�Lf਋�E�<9\�x��/�����G����g4ZK�FPPi��5��R�-lR�~���זeA����ާy�9��|��I����:����l^��Ɂ�$Z����7��1O�	k��ևK��i�j�k4Ϻ�b��P��elw+���٤b�\�Gcԭ>��7��H�E�N_6Y}3�f�P;�mo�s拐+Mg7؛b��'0�vnJ�#�ix�G'z�e��F)��O��N_*(1
F���W�qƫ��]#HBׄղ=������i�+��چ �k�ˉPf9�?\��m��:��5B��������<�L���8��U�<��a��i���h��ZB��H���J�A�9���s�!
'������?�M��$X�	1K�jD��D5�y�_���>��3h��?�s���ib�`�$R�#Y�(ӈ�ͳI�^�z&��^Aa	���ɷs'Zd{�x�7��t�>���\�#��	�:~/k�qD����x�7l{����6�����eu:���0��P�>����!e������Ab�Ymz`�o� ����^��F�D.����#��>��n���E�o��C�y��Z���
�a*aGp�*�:됆^NH�a�_�=%��-���c��_W�2m�KWt&�-��9n[V���seD�M	�Ó�l$%���g=q����@l��J��H�,��8�/�.C��;[�E�D�['���Q��N��DVS�-�l��I���Gf�ʥr/�K��oS�p�&�Q�s?��Jj�))�UiQ���0m�xexj�e����J�y���Ix�%��k�l����(B����Jԥz�|��Ȉ}]e�����&{��T��i^�1������ͅ�v��!�;�_y���E��!�ʙ
����B�����n�J��u�j,8����7�	.��
V�*�^Nϑڅ��hD_�؉�����Q���;>����©>�KtHq�AZlXՂy�հ�u�:]��Ht�i�����g16��h|��f���wvs�)����8����Ky�H��w�S�OA�+�p�m[�		A��+��T)����Qݢ���0�W�� �/n�b�C�v�5�FF	�7G4��j։6��ј�L�-D�u|k�����,γ/�W�I�,�bA�)-ŹR�	o��ؒ���>>.���ɥ��
�*!G���@���
A~�}k�oKK�]"�v��a`�>&�b�]
i�/�|�2@��!�1��i���=��jh00{�6{�x2���e��<��R*��gR�\y{M�ݵ��n80ԑ��U��Q�>�E'�v��Zd_�X'`�G��� z�J���_k��m�lҦ���y�y�l��"��_]cu4�3�#�j}c�d�6��E�C5�֊/� B�1�'!�L�U��s��W�{d�Osg���Q~�o1���~��hZ�W�"^�.�X �rL�oA����>?Yӡ���V�߷G��{�{}I���F4ل;���eP����[�!r^�}?��R�ʢ�S��:�
HPPv����i1k|`Qy&��5h��r�T�V��� Q����p����+<063����e���KF/ �H���#��{t�A���%#����`������qJ7���;���5�Pޝp���X�A��C!�>!�댧+_@G�?z���-�F�o9�� D�t� ��n����M	Ő<0��rr�+�]�.�5~��o�U���?U�2�bЉR 	r��cu؜w��=j��^>�EO�T5�v����u֑rW�j�|�^�G�����E�m��f�(u'���t�>yt���_?���>���U�Y �^������j�%������pV̞S��n�jBb� ��q�ܣ�V����v:�F^r`�� �XG��L�l��/N��ڃ��n�Q�@�ߋ�V[bCs��j�5��(-Ut�E�R�t� p���&�Wuv�����[��q�}�<�����5��"~���ts�v&�o�<���jr����������i�K���vӴRk%1�	E�[͘���W�z�'䪂�'�`�<�	�����EB��/'7s��;^ANY��ڳ�|��]�J���ۉ(_2��6�x��p��T8&�G׼�����������ĒO�[Mm�i<�Y,ExŚBv�ݝ�θ�Ę�1�"��-�.V�c�l�������T���T��dƏ����9��q�{��1����a��Pc6{�/��z깪��f4�&�!�
�N���\j�l��=�)Ky	r��-B���U�D��b������%�&�)��p�|���YGTl�7(���b;�NRY��f�1���_�I9����*�)*��+F��-�ǌ�m�U�=..���4f�f�@<��e����:� ���n�,9�V�H��D�a1��7֗�ۓ�>?� �x]ck�=�ܚ�í��]ۄ:�������i �&HI�#�v���Ѐ��0@f@�!����O_R07��Es�e/HK��J.Gly��ߺL�͙�&T[�k���?5C���Yi�]�8|Z���KqE��B��mN���:F�4<�IXm���<Q�7����f2�C�����Q�i� �}͋��J���,8�)HհG����jyud����}[���&/��S8ǃ�k^<����;r���W:>��<��uYډ�US����&|�m�w�h���R�͕�UY�7)��ӁU�K�³$�(�r8*\re�J'>4*8f~�$�쳒���+�Sw!���c��ܣ�;����.e�:��Wĳ}�z�e�X'�S�����k'�٪=�2��7�n�v�S© ��	�M
PP����[I]㈬@v�T�xOj�(v���KF�m'>�'j���So���<ʊ�������H7Z��}s
���o-,*3��C�<�mq����JO��~y ܫm�ߟ?]ʎ���23�2�:�cAˬ]I8�|��E����/���i��k��:_\K0IpĨ�y'ܾ�镼Mv-�&F�y�|[�gJD���:���-]���i��}��4ƺ�u+�,`?��q�.������|8�O���'�\���^_��ʱo�ps��Ա�%o�m3F���E�]spw�����ޔ�5�^r�C]]�37C�.�w㖒Z7'��9tB}0 x�'Ȋ,�u��٩�Khi��f�f
vc"f�<���;����]*�S&:��L�-$<�$��ܷ0(Mt؍}^�U�+��	;Zk�̲tPL�O�kz�q0�`�&��L)��H3��5q�c'�< }됖>}¶Af��ƥ�L�"�F�\�������6~�����'_]�] l߰x�������9;��fD7ei��dnY'��-�pȑ�WU���D���~�e3��"t�=�~e9iW�促��o�\��yb���l��r��_��z����<J�C���7+
��i����E�$���W�\�ڒî9��0X�)ȇ8�A.Y���&��r��Wp0��1z�:MO��ձ}�����J��;���ێ]K�$���K!�8'����L�b�y��K�|W�%�),�����Q�-��!fC��ae�!��0��e�	zK6.�%0�4,D����j/i:����	�K�qU��0����@N�օ��r�)}�����?D��oF�8}��0;�E�}KrA��)������N/�@�~��ٖeu��b\V$�`�_����Ӵ��{�T����,y������M�	%{ov�ӗC1EA��/��V�Fi1#��n`Bꍹ\*��I���rK-���28H�J�7�������×V�V-�#�
���/U��s�Jpa�����Qb�9�س)k��5@���� �v�%�� Iie���w��YjΜ����=��;�j�Rk�Ty�"��l�~�S�@D~��ɲ')-���*�R���C�B�&�"�)Ȗ�㻝1�YN������r9��9�ǫ��~���=*[���B�KEX��g��ɪ���P��F}El�Er�)�/u�5������m��=��petq� )��t5����d��@s��n�g��,��ӫ�6�N�������+0�!-x.�4:lq���jbh���Ox�B��k�w@��
?��̈́���0��,}<�S�S����@ߌ��ߪ87��=,����~<?�Y�*���C?`<��i��3��)����"Ҧ |�o6*Q�1��y�]�&_6~m|�ٌ�Ͳ[$c&#��F@_�B��Ρ|�j/�h�[�b�u�T��kb׸U��û%PHB Dgk�8��R_r�OmY��V���M��tJ��r�.�E�ׇ}/Ē�R+�%f�wC�� C紐[!*���
��RW�!x{?^[(�����R���π�y>ճ�����'��uS�!QF�מ��$B3�Z#i\�SK������ i�sWl��*��i��z����P������$���&y�q�Ú�%:̙[W��V��5+�� }�-9oHr�����Ye��8�g�֨��[�>vw\���B�w���|�X�ׯ��]��&�%�Z߸7Wʓ@�V������^�[�@�LQ��èEs���/�E��E�������m��b8�u��ǩ�p�[Mb��ꗓ��2]X�);:�����\^Tm8:�"�r4�q��f<#�Ql@;7x �P�z��g�����Z�o>󿢋�Եh!C�B���y��t�o��73��ݵ�֩���+�L�!1�.�E���eHƢ��ˣ�`+�K^���ɢ��Gy��5.�Ƨ��Gx�����������35��:���Il
A]d��}zPoU���@�V�C�X���X׌���,�KAst�֭��̬�q�`Ǔ�Q�8>�?�^E{�B��uhp���}7)Z_��{�4J�S���!R; ���M<��NN>%�)��Z&��;=p�$���]����1%ո����)�꯺�,]��S#\���l&~��S6�������=���ܢ�^�{<���S�Ϸ!d$�mҊ�
��
���H��bӼ	�� x��Pt��h��E��Y����*�ǫ��f[,4;r���QE��5�e6z33���<��i��@k�%�U�����¶22��	��g�p��&7^h�_�pI�Gq<���e��E�Y��$)<8�J+�o��*@z Р�n�Q7��$i�����%��y�S0������A�js*`n.��}NhD͜`�(i9f���T��Fga�Q����{���j�s�e�b�n�0��h.�~���>>�� ^:�U�)��|$f�4X���԰E�F���;�09���y-�7���r�1F���,D���}*(E��í5y��j?
O�J h��mUu����xn,�!�ըv<H|'�/��'=� n����o���F�}�'��gQ�������OK�6�R=�z��p�Z'>^⼢\��'>u��e�m��T�e�Z�4�����0[�w�N~O��{��jC�4B�FC]��Oz��P{��;	uK���������d�X����.)/�]�D��^���5�dMtdN_�M�'ϣ>B��.2��K�o���N{ˠ孼
C׽s"9Q4O�{�s���x;߭F���mAy��c��ݑ����k4U<���`���҇�-��e�ь�t�׬� �XR�J��ʞ�Y�Z�}M�4aT�6KR{�:/� �#X���f��g<�����/��ؘԛ�� �dIli���Hy���:G��-�cy���J��� Aފ!u�J�d�m�+�J�.R{����ÁJ]�L5R��*�0wL<��Y��]wXrk�Pf����WW{ݞ��ێ	�]q/(Ģ#翇���������.�`�ˇr��4H�y�tŻ��Fj���eT�:�\���.n��_�u��-5�0�Y�:����QJ� �-� cލar�?��ʡ�)���)g��%V�wa���)�mi�ew<F(�������ndΠ�Ӻ�T��>�
򽆘̫�D'&(#f9y>�X�wh��TF<+�J?a���?Q��5�d+ �A�ɢĮ�]5�ٺ�j��OJkY���w���"A8E���3�(yF/ݾ(_p` 0hr� Iq&j'[(G�ϱ0.MV�/�	�#�h�)��]f ��K�HH��")�l�p��<Z����\}�:�3ͤ������7�43}��E(�Ո#��8�Y��"�����{�]0��ق��}�u0l�ہƻX�T��K�*��Z�<Qi��(��Ê��J��+��}V�ڣ�۶a&�JMd�Y�_��	��f�h)M��ҸG����I4�TD�f��V��?JU[�\�N?���Y�ᕄ�w
���b��fZ�sW�#����)����׻{�1ܣ��Q��At+�Kq��|��E�x��y���4"�#MT'W��3�~]�b�1��v�j��Mٙ�s4��vh�Y"�8SuXv`)��Ci�CV��e���x����Q���1u��!����>����
�xV�^���`���	�P��\ߥ��Y�P���=��K;JA�|�Z���	�o�����b������Տ�ȉ�N�r�=�)i��1���ڐ�Q`��&��U��cK����'�M��0������2Hix�(�=\e>E�d��Fw?����M/������q�x���4o�xAc_G��[���h�zȩ�m�N���zM��2U�R���YQ�,�U�OjA�ѥ��_��`��(����L�/�y�2�����`�� ���^���c�<۶�"�!�a�ų��t�S�
K��U����E� �@�����t��[�9"e�k��)SOu'�]����?J<����^���DSJ+|���[�1�'�(��\�d0A�p��*:(�!da�V���$2Ak�/Ҵ���@!�"%>�o��<SR0]�T��*k�s�u.�L��W�}IB���&��b�c�X
��3$�
�����/t.�0����5�`D׃G�P��b���<�Ɛ�S4���W_
�IF/h���m�xDܒ�݈�h@��ʵ�VF��|����Μ����s��[��
�{��" �qM�ε�����)V�/��[$��д�j$�~�~��m��,���0A� K�$^��N5S\�O4E<��FIH�䎦�U�/W�g�Iw�F��|��0������x84/��"@��Dߏ���w>���@`r�Xv2�Ud{e�Z[��oB�� ��>�ec��y�3*rCX�8����t�_����Pӳ�7��;�#���K#Z���UH�JU�d�9ڍ��8<��m?�5�·9���9���B�;��|��X�˨10�TL���cY�)�B�� b���g\��B
�E���`z��f���fEy�>�q&(+���f�/.W�E��o�fv
���M�)^	�;�=z�Ɉ��d�l�#u���?�b�"�"���*�Kjr�
&�0����u4:���e]}��]%��wɐ��~5�I��+_���:���8�V��N�.��4|=�b:D���uAZ;��l�+H�s�0*k�ff�|E��bs�1�2��5!�4������3D::ի4��U��\�a4�����..�pd:@ mK�6�i9�y�Z�si�jd%��8�{�V�P��a!E�j����l\�m#�.* �j�cht�J��[�8��%���o�wq����ݾ���4�A�H�	��nO8p���(ne-6�xSn�Wi��i��"tߊԗ#��?R��z���.�t>$�\5n�CqnW�%�xfj�]��6^tF��Bc��Th:�t;}c�+�f�g����o��+>�歭�e�i���`��8�-�@�w̗�!B���8��@J@���̹9Xh4�,?�'&�u��	hx���/ɓ���n��n�u�N$�.��p���&�Ŭ�GH\���]ݏ-'^1��1$l���6X�c� �"��C&���$ƥ�؇;7S�eY܃7t&�o�����	r������@����e��iQĬ69��Hj{�8�D:����A�ؿ�U����G�;h��F_����C�&Ҹ�>��yٰ6I�a���ޚi}�	��j��:�4��n[W(�l��>8��#�����
�0٘cf�6�zOj�������מ���8<�z!]��+��I�=�y�*A<2J9��E��n(�m���s�+���(�Đ��-���_��V���m�A��m��L�+�6�}O1E��m�}jR������Ư]W��~��ts���^eG��m<�J,��P�0d����	�r�t���g�Í���Aɭ��4�/����N~�"�!�Xr5e/��B�iL\e�{o�v����������o��էR&l�\�*	����T���6g5w!a:�E��(٧���)H~88��`�?��E�Tn�u���N�k۴Rlp�L�r����L����w��A�j�fW�<9T�Jl�B�e��F�f���i�*�j
�����b����=([�a؀\"�˄2�Ov�7��e�s"� )�kԘ�VS{<l���c�%����k�-~<� ��rC	���o�#��w0Yxr��tvV��(���:W/5�ֽ�}
M�I�3�z�َ��W�

K�H�_g]	�Y��c6i�v����Y��En�֩��.c���r1k��ִ;Wa�(GW�vF����e���0�B �W�D��V>���}t��%^���n�u��n�'+�O��o�h^\�I��w������Y��v#�"8=_����q8�3��]����y7ca��������^�t-?Ƚ����� �e�g�no­7�%�H/�C�)nS:`���M(Ҋa4b�&}�A�/�z�\ɢ�� �:f/��I�3(s뎩����nP��Ú���2��(��Pg�=I��?X�#l1{�~�C�%��,���''����'�Mk�	U��h�Bѐ.���3�%EӓbC`��n�.�g��`~�V:��M��s',e�(��yT�C �?w뀘X]@kޣ�#��ܵ]�qN��m�A�<��Y�}�r۴��� ��6�Dx� �䬀n��7����K�YI�)_y��o�Kq�⼲�	Aq1��Hg�	ȋ���B�<�܆���*��n�J|�꿡��"`�������B�6ڪ�bպ��ť����W��[5�d��TK��`�[�Hp+w9
E�iس�������z��ϝ1��,����D��>�j����w��ڒ M�8q�zvy��`��n/�/�ZfJlz�1�d�_����11̳�O�uƹa����:W���jZ�Js���.�(l-qs?�΋Go������E�K0w�:ᣵ쁖8=�;��	�܌�ws��G��U����%Pi��0}6�����T�$P�Ơ�Ķ)9�N{����a��h��is�%��-��4��ʔ�Zm�����s^�����J�k���#��i�t� �o��B�;)����z��׼���raj-,6:A	w���2}%y3�" jU�k�t�#9�̹� y$T��\�.f��D�̦�e^6p���ј����wd�� Г0�^���j��r�=|[ɱ�w��`��0)<��t)�\D�����B�W=TB��}&��"�fY�K�-���8
�!F�9�u>I/�I�=����i\�7��a������������jN*z.,�1>c�y��� ;�.��<�w:,I?��s�7�LH"��[�ǀV�1�#�L�_J���}�[g�g�J�? ���k;0�@n��2���%��)�e�5;�u���&m���]��c!�c.�-&̂aL�9���5���ȰI�,u>#�)�lgI��i�JKZ}}/iOl�8&\�CQZ��xՂ�J����)�|z���H��[n������$����+e`;;���A�s *|�!����P�*��UD���	�	8��C1�c���\�i(�����a�>�������JT*�=mƪ��%�I5�i@g�FF��e|O	4R��a��w�Uhx����'V-�HU��;u�R�i&߯]MO����pg�!�8�?���=�ԅ^�4,������D����)���� ���)�(�ܝs�m丐꒕4�!�9���T�,�LN�ㇰ`�PKOMt��D��{�+����p��v7��/���6����v��������ZzK�ޏ`Iz�۩-��8H ����X�%�[�8�������Xq*ٚ�=T8��z]6�JLE��~�E���L����3��"���N��s=�"�J�=7<X�~Ph��g���1����l5E]5'D7�����:ޠ� �"�����]��������J�{]Ӛ�ă
�~_Oĸܠ�4�(��]"�a0��VZXs�r�ծl�80�r���WQ3@�ct�E	�"�i���� �A#e��Q�π�.T_�n�\��l��F�W"�5J��[�6P�� �0���>�3��!��|�,�S��e/�KjMX���6?Fbf��ڌަ��7�ѥᶕK�:}�[��V�ܒQ�Y�<Q��_/�G�Rni�(�<�O��(�ɜR}���-�r��҅T�ht��D3�a���i�K=�B������������(ẗ�{�p�F%=��`����VH��p�cy�K��\~û�/uh�Fwk��cT��#Kk$�R���(���>����Z|ui:ݮW�c�)��G|F����hH�F>���G��+�'?���%L�S���8�u���٨.u$�o��c���#%�(9l^�V������z".i>�5�x�����s�����;M��0+|����[+`{��An����Fc7X��t�0k
(�!��H�Bø���l��v-�ފ�T7>�N�wE�iM�釸��L1��8�@��] %�[�P�������Z#������a�"�
��D&U�VE�jּ	6�Д5Ml����]����g�D�p��K��[��b�:9w� �)��щi�<������C�X��#�5- ���mN���<��gs�9���/!f�:H�3��y�
��L	sp��s��2RY�Ȓj�3��O�_-�� ��=Ȓ%'+�4��|Oh�z~�@��`�P.���S���Yc�CI�+���]\\�ך���G��u=��Y�E}��n���b�6�7s�l�+ٳ?��	PRU���13��e�Kd������ne�)��%D4�B�Ip��V�L�đQ}�&�Q��(ﳃA=4<�4�0{��q)�r��uzt�d��(��[ߏL,п\/��X���b<`�r�y��=!~7s"�5Mr�E�,��#,ɤ4&��Y�P�"���^8�Q;\.�,�mR�@����܁��XL$%�^��>����z�%�cD�`	b�Y�LdB��У���]ο���� Hk�s�⚙��JT�EfT�������{jk�,�/W���3)��R�^��W�:-W�^d�v�:�z�̬�lя��ѫ��m��R���؄{m�5`�����à=l$��W(����N���Q�j&׈@9�_�D��̵�#�xm؍���+�=��Q� ���x�!�=��{^��FSc��`OjY�D��,m4*��V:~�vI_�4�K}�Z>���_}�����X�sb	 �h3��n�P��|�I�l1�g�?���-��,��~b����UB`��|*B�r�S�	�P�{�����1gV ���J�xtȻz��c��ώ�-�����B��'��wU�f���9-Y�-�`Y1�ŁH����-��s��E�x35�E��ePvJ���S�-�����,4�T��HU��P��a���U�v�o���h_%����aK��|{�&{�x�>�d�׬�/��l}�C��P}��p����B��	� ,�6x�����\̻n0"¢�31��fqg_��8,1�,e"�S��r�.Q�"�3�2��UV�H��6|E֮�y���ח��W��$�F)��M��<_�xnf����j �ۄ_�hZ���?�sc�(B�/�qħGd�����׀����WE�T�
�bI'�hM��4���b����K�H1"�ڪ�q{CO>l�Ōk�C���^��oP�5�X)hHq��)���^�Ġ0�ƍ0�U�1����_%5�oJ>KT�{�p'�9/�G:�Wh�*Qꥩg�b�7O!�f|W���,��)��j�����V&��@|K�/@)%4����m�د����x�)��U��g[�����C	օ���!L�ɸ'���B��32��%������mL}�	(]ުAh�^�uSf�vٙ	�9�$(2ݭle� �)�J�3����W����H.�"�<�({c���B��g�߉�D�t�|QQ�ٞ�BX.k�`�x4Bo�mJbcI�BK4�|N���y��m����Z*�Qo�Y�����k��M�~�V����6�e�h`����2�w��wLd�݉�V�	dq����]�HX�����#��eq��[iAi^:��se����m�;6&v��٪sj���[P�9���}u���r*[tl�Y{�I:����n��_;g/�|(�7( ?OH�G�Is;�0!�y	{�J�$0��r�]f�B͖����0��v�'	�{����@���!����Y$"�"
���n�V�z��zox�U1#�����"0^R��=���ɇ�EI������7b̕z�W��5}�ws�e��W�--�vI�g��^���[��L*��؅b����x�.;�h�f���Җ����&�/c��B�,���R�]�Ѱ���w�gX�>��x�c<�Nr�[�?ξ��k^�B������/A�B{��`J�M0���Ѣ��1C���j��E�X�׷�A��^�|��{ֲA����D�8�����=��P�������_�wڶ�(
O��ƈ+K�^��v��=g8�e_ˠ,Yh�g��ր'�&X�z����K�߰�X�)r'S#mrI��$�ÏQW<z�C��9d�AC^�*oһ��(9�fKN8��^��qq`��H�?n�y�y�c1�`A��/kF'ԟ@\t�4}�%��h�"�Yl��8@�`�T:��v.%�z�G�yU��������ע��lZ��Js	lq�Lq�ַ��N8�y~͇gB���C�B�7hzٍ�i
Smar_kΓ�$�Y��b�׿yW�����E����TMZ��#��T����;�n��QFj�C�J`����xe�i�g�*����k�8��B���$��>��G �����碚����E����ܒͪq��nv��C�+�x��>�r@S��QJM�I�;-R:��]����[�]�Ru���>|jюs9wIA�"��~@ڂx�^��J�7�*��!p��� �Mlz��ը:Ç�����)�KF�r<�>1^	�Jq�ӟ�ko��Q��q$Rc�]��+���K	n[]z��Y��a��ʐ+� ��w�Cg��f%����Wt\��.��K�]y�>����@+�ɑ`�6�i��d��;�w�J%�u~�x�Uh�%iz+�{�O�s��cY�5M>�M��ӼW���c�K2?b:�(�͞1�������q�ٍ���
G�.=ooV�b�g��l���&5��je ��\�_N:
[����`���,9)�j �!�ď������!�=xn�xXp%��O�j��:?�W [�G>X�f�Q��b�.L��l��5js?���@Za"�����B!�(���uɧ�ߗ+h�~�J��Pp�"��fE+\N�s���K(찣5\���xE�]ΰ}���
�k��q��G�}R�zeKt���݋�b�?Kd���p�D0i�j��R*�(&(�=����D>,��GH�J�ۍ�p�F����ι����	���I���ߪX�d�h�6h�V�����:�|K��y5r�*R�;i�mY8c�e�2e�u+����W-�X�ҋ�<�=X�A�;�K-��].�5T\p�OW�:=�I�%��{��_��ǝ
/��CR<.idhU���i�&AR7����O��o3�C���-���C>�R2��o�ڦ�9.LQH��y�m�*���@��$�� ��*4�UM� P��G���(LH�H��)V�U�ķ :k�&G���
z3�W@i�%�	���b���o��(Hﷳ�e8E�2���@fIjB�߮��t��b�P���%$�~� g�t�@?�8GYG��v��\�<�D]�P̽~)��}~��~`�J|�������u9�}L^N��\��^!~*f��w\���JY<u��Rg��KF,�>F�ˠ8���3��M���S�����O���GXB��t�%bBP˵�(�O5	�GE0JeD��H~�F��&�ZU��"4^�p`����bś����V<ۉ�-����/��!�?Ȣ�E�]w�M���5aty��<�p,��l�'?;ij�5���LX�6�>:L>O����-v� ����z��jm���P�J�(��7	�����*���3r�+iw#���NuL�;W�b�ֿ9��av��~�����Ůc�o�r�������p3��φҍ(�;�k�6�.�1���|�eQɹ���W�mxlM�T��dtߒd#���=����]f��������&�6��*���>�����q����� W�A��tap3]�J�e��l�rQ����f�����/�f�UX��x�^�]V\Q�!�$e����r�/8�	����E���ac�g��xZܴ8{�BpѾ����͢����T}6�n��TJ�v�]-�A�lA����-�L��8xk��ퟣgH8�Tz�0(Qž�_��9(~g+�c�=F�׶B��l�Y��l��ͣ���@a_�	����8����Y˶/��g,\�g1��F*^�G>�~>����
�=��5�M+`N��7�����\��c2�%:]�T�W��a������|4�6fvy�3�:�=��q)#3GOsY3\�ߗZw(�*r�;\���e�J��abQϑ�9����q�%rcZ�}�h[>4�K�|�Ac�f�gJaY\�[9����S�e�c��Y͕��"4�� ��g>F���Wܕ,DZy�3��� ˿�s
	�}�6�йB	Cdg$���\�3	�m_�"iS��7.��ꊜ_ځ\��5I��J;�L����Q��4���Q}n۔��J�$����������(���^�g��љB��y����i�/*���Q��H�R�,��˲M�'�V*�cnN����\N����%e�_��I_���/!O(J�r	Z\ނ��N�7"�u߉9R�ʻ�PP���H@�	u�3n�}b�˳!0�ݒ�A �8XS�:��?�ƴZh���Hy�K2�U�������E���+��bh쒴q�h�*�$D����2_�� �)-��Jްi�6�U�to6�����G%q��rg���J��?��2n�d3�-~;ئ��1MQ��c�kʌm-�V.�t4d��o�JW�Eh4`���^���Ͳ�����h1#���?����5*$�x{j��"����%k���ڄF�iT2�m��aК��l��r"�S$T��A�/7l���8=���s7Q�r�r3b���#!=һ���X�
E3݆0�UF,��ȀpƝ�f��ɖ%��>��I�luqu�p�/g���
�����6sd�h�L$��z�a���������k���ȏ���{Q�����q� ��̵C��5}��$apI3��Θ�)�R����*�u _�sgg�i���W�7�;ظ��vKں��	 �C�T�5hy+.�t�R�g�C�9g̴n�56���YU0����������;�����JD
�f��WDd�ݰ�����g�J4i����_}!��;��^�uT��Ѿ�����v�u�0ȇ��7�Yл��xONl!�̄�|M�%5�޵�͏H����I���3�K1�DOZ/�:ǒN�۟�H;��>>��}��Ԝ���F�G�@��^]Z�䵂gB���#`�+��M�?���eP[�����`#{��~g����Ƭ���[���dG+�.3l��8�?12�X�7y�l��+7j���Y���z�4vfrYܠ��$@�u^����cB�5!c�pHc����r��&�45�w��h�v:;�5�0��32I���d�,��v7U-nQ��2$�6S��a'a�M���.���ʊ;����g��|*<j��QC��꽌tLz>���G��?ы�M}3=��6��r��+��GЏ�B.7����^���T}�7�����H��u����؍/غ�� Q�ܵ0 ��-�Mw�̜j��w���%����mSG]7"�.�7�|�RG��$=a�Dd7�Al���jik����5Z��^17��W�s�����/8X
��=�Z���PI;�F@��y�Ͼ9O�-��"@h����FU7H5��`0���-�����2�:�D*U�i*>�Cf|)Q̝B�G��a�����K ;g��l�������k�ƙ�=��G�PJ8�Q_ �����ֳ��B)�(���]?0DI3d��)�U�L��9��ϏJ<t+�[::�hg�6C����.q ������EhR���TfgʤQ:��u�3��\��^�D}<ڈ��?둃V;�g�����:�i�^R3�x�iš�K��͓d��ɜD���(|�|V������: ��P0fs4մYb�Ny����e��?�{���x0� �g�%�����x�Y?����A���e]+��^$rd����������oV a�^j�5|fD������Eն�Aַ�?:Z���&m�ڰ��΍�pyT�)�Ǔ���:�/5�%9z�F��(py��;�����<�/B����Y9Z)��9����эL���e�~����#b2Lbp��O4�I�ٲ9��{���>Md�D$�hL��&�ҝz�iD�X����1P�M�w}Ðq�E��Dſ��)��]���$ڧ`�y�����FR-$����k`N]-d����{Ş��,ŉ���0�1ي���쀠,L����"����tybA��1��0�����T)r^��l<V�iwg� ��K��Bed��HP��p�{%���Zm�e|�E�Z&��u�@1\	�R�,��F-ױD�Y�y7J�u��RQ��.��w\����x1�T`u�2�s{�K��f
nuZ������u^A��FU���C���i����f�$A��Z`�a�S�H� ʎ���8z_L³ �Jɐ�Cb�q��g��ٙ�_��M*}��y���b�<.�Y㐯B��s9-�g(�{�{}�[<�`��Ma��6L�J��4c5�g��۽ ��!���Qy�_j~ ���?+zV�'�Y�B����4�I{��'.J�\gDı�������}��"����h����8�hp��u�C����n��O%�1Ԧ�j�v�i��统�.��r���������wì���bB���!���ӥ���X�gTُ��#�F�xHӁ%خ2#>��MY���'  ]ޝO!X��q*�),_e��ʙ�5�@Yi�+��=�)5p��r �JOl��`�a�ܖ��ݜk�W��SG�=�g�!�d���r*'�.Cg��7����.u��"h|��qfr��ۑn�`��C����=����Wه��z�Р���`6i�4M�����>(�Y���@
C��C�`�B����cu������9����M���{[�FCb}m�\���$ܮ� �e��|���f�~˝�j����ūE�<m'��9ۇ���߿���K��-���:�C��ځj(m�Nz�ӪK�.S�c<j��2�`zu� `s~kC����q°��oPY`<ŷ�VG����;>�
YL�d,���8�]��� -l��� �TN'��m�f<�. ���Zz�Ŏee�=��#���9�*��$��r��b����#��������B�D�#?T�7g�Q�=�E�ֳ���כ;����/��Z�@eUgo�2ٵ�:J1ߛ\*$\�m;�|^���GbGq�G{w�X���C���xv��	d��A�?ʟhf�6�@>�.A3wp �]dl���@B �h=�K�&8!����t1)�K�j�n���X�<CxX�~���<�ˇv���F%���f��e���Eӳ�8x½�C�iXa�Ԛ���'�q���S
TԬ�I�R��;�䡟,�ca78|����ۢC�gc�7d�X�1#���:�M޴��]�|�,�*<Rd湗Qj��wB����j�f� �֥`�}���0!�t�)�瘗N��0��6W<���WI���y�iGD��Lp�Gbв�rex�֞ğB���>?%�H�?`��yT����W�_��Hr~��T���_�"���[[�$���"������ϋW�<Rٯs��?��'(�kz[��S2B�DZo0ĵ����{�i�'�\�е���Zg��&.�vQ9_|��;�~o�p9d�r	����Z�텛ci�QO�Ŋ2������Ҙ��Y>������7�O
>rdC�Ⱦj&�oN��F�����.����/�2�Qf�ȩ��G��&�b�n;���O��W�t�`o�)��S�:@�������Z=n�e5]�H�s�N��c�k�b �2Cb���8 {�����<8��&�:"���]�|���5��V�*E~��Q}ve��\ۜO�t��!��Z�M��L��#1�s\^Ы�t�
�tR\�}Iޢ��^��Z����y���qb"p���W>̢:)�I�ϋ$�����e�768��(�I"�:�0�N��f#�<�B'�Ƈ_������� �v�p��r�Ɔ��ig�a9@�f�7gwu��$7欯���_c8�8Q飺={�%�2Kc����@��_�6��}K�O�5���x�0�d���;�[F|tS�w�t��E�����'%aA�(�&2�w���
�ʐ��\�e�$ے����X*������"��1�:d.�,0���i��k�@��n�y��<I�<� ���4A�~�'5���م�7���0$]�(�c�������՚�<�p?j�F�"gj����=��V����� �"��j>.ɧ���I��
��ACm;Q��ǻ�|2!�97�uC>��Tv�N�[�v�Ub�����M�@9���xۦ4w��nX���m�v,ZX�RV�Y�m�v��]���R�,��}Yn��7�����i���} bc�������������Z��_����wQ��N޺�����8��M�k�+���=�m��-Β���v���5�2����@*���~��*~xUY셞n�3X��[Sq�^~�uI���8oШ�-ۘ��G�6�M΋���l?'����~bLJ`)�^�.�A2�mg�a	U�Lݽ�GT�MOd9��}�ud�Ne�����;3�L��K�!�om�.�b{k-�t�x�� ����f&6��BQ���eL�����z�g'�ؗZ���e8����;�< 1|���=C���YH�jV���GY��B4Ux�kg]��B!t��wV8/+���7JOq5!w�"�[w�� `|ɾYX��d���\A�c�,o���f���OV�l�����r� ��������ʯ..rbj�d7qMC�,���n#�g�>\�x8,��L��NY��>ġ�|<#� �4�V������J&�Ҩ���T"���2�0��*!����)Y��{>��>�qI"o�>�h;�������ī��:N��d����!r�s�Y)<!���|�J"�6ĸBߓ�X��Α˵]JS��Ԅ$�G��$0�_�!��nP/z�=cz�D�*��R�Yi�{x�7
�콆Z:]�H�reW+���,���.~�+7#�c.a�Dc��Z�}+� '�`����Z��S/41"ԥæ��tQj����d���s�#�m$o�gr�.�V�qe��7n��l�>���c����e�R`P@:[��<����$��mD`�-]�޼$�If���G^c�NB����2I��:rM�9s:��'�]�l�k��G�����"W�`�$�7��[V�6� �ϽMe�@Ԧ`뼸y�৹`��Ơ�Z`Њ	��NL{���r0��܃Q�*:�s5�t �(����u���`��V�D>��;��u�$G���c�U�өA`��9h~�\ɇ��6���X,��H��s�ھK�̐�"� &��NQ'� K4�(O��bWo�����E���ȱؑ?�Q\<�O�+�6j�5���x3�]0����{�|Ƴf+υF�1���^ڭ�/�ft��򞪕/6�l,�w�������h�嘆�P*p��g+a��y��ɲ��1[0�:��s�u��@�d�D��-�/2g_W�߷��+|�"�C"�*
�]���W7,�
��Ϥ�S_�yJ�_��.�k�qR*�!�-��ٛ�QWĪ*���;Q�=/�(��؜X8|��桼�L,�&�|W��>=+ʀ�fh�|>�r������[���{G�A�r�Y�-�z�:,:�b?ӝG������ �4P��:$�i���t���3���C\�n\.��$�j�@�$m�L]9Ę�P�Q��a�{n���R0$�/ŖK�/m�U�B� �Q����5�c>��n�	��'�EtP�VK��f��D�<Bu��L��@fsk��v:&F�w�J���ԩ��S�g������8�X����Y}/��
���_ݱ~b�}�L	�;˭�����U_L5�da]������~�-j�OSu�P1c�����5~��x�U�����tî��㱔�0�x���h��Y�<���\��R��$F�h���}���%'�ን���1;���;���,%��d�X��V�;p��8�{`׆`K�	݅o&�\���}v�}�{�;D�.*��%��#5X�ysk��X���j.�_��D�d��|�3��/���١%z��-��HB�^�b��o?��SyS���ڷy���%�_SH�D�*?r����J�!@��J�bp��q���R�bzI��^�{����g�\����Ԭ)5#�[c����Q�t�S��5�S�kF�jY�.����� m��&M%?��Ek�R�R4�r�z�&�#�Q����ZY��H�`܋������W�H*��l�xu^�q�rD��",��3/rr��ǖҞ��Ɠ�p�7b�YA�y��8�o������#]P�#"�-y���v:��%v� P��9?#5�vf�7L��\�пZ-����<��/V��Fk5����7PH��v�O�+�ܝ�%��A�x�aF����!p���40��z��2I�'z�x3�C�!�(c>�x���Kk�$�*�*�Z��NҼ��HҢVa������QO ��JGOdG��S�����������{���&D6f�M
��̤1Ysrh��\8�@�/�x	�J��uZb������|Ŋ�+7�9D��+6@#:2��Bܚ�\XS�'�O;�` Ν��g���H��Y��)bxjڨ��O45wi�y��y�o���)��A�!=,�<�H�5@N.0Iw�2�a"#j�(�o��\Ɏ�����M�w����4&��L�V�A����r�⭺������������Z$���Y=��a"�jR(V����Z:rbh�KsB]]#���!F	��H�gpם�����EFiH�ƹ�a[/���D�;��%yw��k�Z�9-��f���L�pO��𦐴��5���h���塛0�n������"w��	h]��-�n�C�F`勞���h�.t�j�B1�9�5�� �h���4〜s<��_lV��H��J��3DHh]:Q��zغ��wn��4`)Rvޗ�XW�+�,ik�Ş�I������N� QC����=�É�i{v��dF�ǿ[''@�gGy׸W�����C�Hp 9db�s������ L��D�2H��QJ�}������ ��=AD[��Ȏ� 	8Ī���/˶�� p���9ۙ��xρ�3�O̻Wk5 ���|:<^�� ӘH@:G�M�*�f�EWq��q>��W���s���KǠ�Ϻ�	���%�3����MjΧ-t�	�ĉ;.�W�zAx8vQ�r@.�\}�"�t���`*��ք*f����L�T�Wl����;�����5Ra'���~�aj[�\}"k��C��N*#(��w� �k�rL7���of��z�u6-���	��CW���������É�c�}5p?!H�����o�Z5����PJ"�&�6Q)	�:(a��ʣR�d7����^�%�ah#����a?��� #��_�$���R)�ѝ���=B)�eNƳ���~0���6Yӟ�7��M$���|]�%�l�7;�:�ڋёU��(��P2��������Q�h��:���lOH>2�����-�9��ǚ��ԙ.�'�Z�ޫ���_Ңie3Bz){Ս	ٯ���\<qe�q "߃|�_2+x	VeȽ\��s�X���@�;�^��ϣ}�:���gt�":���ߌ�]R7y@���{�A��w�+���QR��;y0��I�{��W�o�`��F��D�! )���+�{p*����o$.h(q��"ז1��`� �V�F������IE	�ֶ�xu8k`3�ĚC�e=����H�{�t%È�/�6�~4�l#��� "pX��%-���`9���&veN�<�^��;>�G��s���G����7���X������5��itn�mvV�{��Î9�����K�K�����
6?���r(�婻`#3�����]]g`�X%C�-/�A.����vb���C����ց��+U?�v�-�U� g'�˵P�����0�{*��>��=<�UOpE�
�����!yw u6��ۚA�?�`��k*�;��`2�u�{���,�ǻ�����t���iϕ�$"���c=�惝NKڡ#�4N8W����[f��WB�	�`<.rM0��$;�����Td�Ѿ5�����dr��!��tW�㶓�6ŭ��m���6�]
�GEAt"����,s�����W�QP+�.Z
����hE�ZU�7��	���VhA?���5f�Fx����ʝ*���b�Х�*ܽ�Jy�P��D�\��'�����8�7�go&��rH*����A�<�����IK$�, ��`���5X$�Ё�q"���!��g;� +#��մ���ڈH�L�z�HP*�����SWUM��w#��"�[މ2��yN�Ν��]�赗`�w����F}PwЉ���y�+�P*��!�W��G�E٦9�_�gUP�Z���B{�4EZ�^{	�`�D=�8�ZS[�WGV����dP���i�z�z�3��/s��$��ƌL�G@��w��} ���m��e����q
_8i�H����j'콢�~N��r��R�6����d��M��|Y�B@���>��왨�#�����}�~6n1�C���m7mR6�@zꙅ[M�F��`ʘ[D�6
�+k�k���~$���h��L�*�rihF}���
�a���#����Q�pU�5�_[p7�H;��L�-��D"%\�)%0,�Uޥn�	m����Z�eP��\� ٪���i�4w*�rA=��:�+:L��m$�TS�{G��������h
�$>��|���믾-R�=<;�zR��0.:!��uK�������jT��:`�.m�nh���B?��ib�uD���|��)��G nD[�RŸ&qhNr2D���CU���lO�' J��o���܇���#B�(/����7ba�Ʊ!g(PՓ#�;OBk貽���%L�p��>$G��P/	qh}9��г���n�]��梌�|1`p���)$>�b�6��~`��!}�D�O���i�����V��O�p��r���AOGʃ�"rI��C9fRWZ�X� /ʻ���ۦ��zw����?�k�����} w@���E�ɱa8�1���䡖N43���>G1�QE#�SJ-�<nc�x��=��X#�aT-C9�
���:����k\M{n�A��ݬh��E�~M�sX�B �	iD݌q߻���n�5������򞣇��E�$����%d��O$���{�
��Ѿp��J��������q��=��wp����W���z`����c|��T� ��,ÁD�Q�j����ͧ��<�SOp��G�%�p=�nY�t�!b�ܘR�\��MR8-�N��/-+�����k�>M���T񌈨�嘦�Uۗ_�evH��R	��z�v'�����Ȗ�i�_!m:���b��L8�#��n�l"t��hLHVl�^*�˧ʴ�da�^PQ6B3)Y�1���m���}~��"a����<� �q��sM�D�/\�f�b8^be�s����y�Ž�!�z�ng`
�\mU��RЄ�RQk9'p&��H�E#�����p�j�r7�C��g�B������f���;��1�6���%�61N(럎�f>�$�E�V\�Ǘ���p���dbv�^�L)�N0���xmGѓ��¦�9�"�%;}n������&��.��d��V8��'�,��BwE.����L�R�s�N����p!�p+�C�3�{�nI�'d}7���k+(-����{Y��L�,���-I�3f7H8SD^$zۣ��P2{��g�()�Ԅ1;ڲ
ӳ��Eyԡ�9���Vx��i1�+m��� y��I+L��=	3�C?d�~ɍ�brG���I;��&��o5�� ��A9�8F#�v�7u�Fn�e8�Ġl� ]s�y�4R��]�'�1Q�k�E t��V\R��V���v�]��?�8��	��_
��ⶥ�CE���\�jO�{�!q_ߓ_ʁb�H�n�$��5���0��9��`4D��;�c�zkZ��I����K6��r惨"�?�mF{����..��;��PAr%�|���ӡ�+�<�E�w4;#ɫ°4�9������b"��($Hu����.k$`��K������е$��h�����jOg ����<XF`u)�Gק�H62�B���BηA����L��|�������/~���g�wA� n!������Q�AĀk��;pi�D�oz<��$>���;�ޮ\��Xj�u������2Z���}�M8�th�U��j,UH:^����.)�%���M��Zm���r��ez|�Z�=V�ͯ��bp�T]W���%���E��(ųtM��i�L4�d���t���f@0���'{XM�X�c-�U�TM|J	�H�N9/�ea��"�Y��/����?|�u�+7�@۱u�J���I>��c�y���`���3:�d�@�c��o��Q�F�e���%G0���0�����{����Cu��?>�^�چ��G�+��ք$�+i��U��	�`4���xO;@q��	U��gʫ�������7�>�2��<\yExZe��/@J��Y���^����u��Nܗ�/f����d��j�%r8~S�$�蕗��;͡u���7�旑�g|���,�G���C֠��y&>�����d*(뀳����1�zFG�����J���9��<}�$���B���.��q����z��HBE����ӈV�����?�b���ªƶ0���^^D�k���p���3=��~�\�+;�b�b�9o4�Om�@��0���ͤC��+�VYMi�����BeMR�]�0Q#-���gb���ͰED�x&�+=q%�Wc�p��L��u!R{��S�v�/��ˎ��z�a�"Dġ��`1'
�X�c�.�Kc�~�5h	zX�� ޺,H�qɬ���B�� �������D���Z8K	`<�9?/����V���Ev�\*���������+0h��o�F���ͦ�L���f��V5��:�}��M��"��z����8N�l�1��6:��O(.~�&l�ySY�<�����a�+y�M	�As�8�*��ud����Cqmw ���6+ߡ���n8i��38��wq��W]`�+�H��}���.N�Ĕ�1-��.�	��Q�qd�j��Bj
��;v�Bw͍����fVt�z�Hx˶�R�ef~��EK|�	,�8�3��X�bXF50]�Ld��3bA������dy� ���O���
���9J ����R͉��J`:�x��!�y�
#*��1�j	��r?>!}}[l�\�\m��K��3a��?m�r}�Q]�%ފ�N�ǖ]�U e5E	i�q�� v�3�V�wτ�+E�ɵym�:ݚ�u���P�x9]���Pa8Q����%�`�JR��3,��SaE�2��!�����A��_>��h��.��H�Y,[��e�ߜ@�#VaC���ɠ�FZU�]Y_+��עߡ!j����Ѥ���m�B���l�.�x��ޛ� ����c���̪<����:����k��u�G�l\�5� /���w}Kв@��F�Bc�rg���>��F[i�=i;��g��#Rp���{�C;qB8�ƿ�(`��w����F\z\��7���#�L�J�IR��i B��`�j���c��f]���ޯ1\�.ѐ�^�p9/{����;�`r��B�P�x�ۜ��W@b dψ� 'f�P�<g�&`�
)�UR ��A��7��1�#1U�+sq�#yS}B�FK���*��A�8r�~�bGQ]���i<�##lX��)�p�!���H�;�4D��wt�2=�d��N���_9-r�`�;[�����h��If�	�� �^ھ-�NH�����
�S�E�ֺ�Q)	{r#I�[�Hn�O��y�����%�3�s�U�C)cC�� �Q��sw�mw�Q,J�e�x�IƉ>�poR��2�E�ݍ�A6����n��H�2��hNE��w�J�ر}�	�Y�GN��*�=Q�^%�}C�-����%Jv⊪H���={���.�N?�UE�dK��b.�V��dS`ko{��!��'�x�¸)�H��8��f0mv!���d�<��_��e��*|�^��z-����]C/�����1�'��4b�ӹHd�Ț��ת�Ai�5�0��*1B[=�v	�)n#ڴ_���"x��2�'/�^_K[�qr�-�9.iXG5���m�w�/^t6��^&h3��3��?3#ߟ�K,+ݗ���	,duФ��5B
ג&���@b�ד;���۲��(�c��n;,x7Hv8{����h���Ib����EW>8�g|8��۶� WL��3�ۃTM��S���;of��&�Yph�nb�H�}��`�kG�="kiRqt��ێ�L^��TN�!mשQK���c0��?W�K��r�,��T�P��5��#�ĥbn�9J5�s�V<0|u��eL��7�_���Ԝ+���IzFd�����h��O�����X2h���O1���J*0���!�oq1��֭�QSR%��y���h$0}��@Y+IW��۩sP-�il���<f�"+�p��ߘ�4R×�'�T����ʲ3n��`� ��a O.�>E	�Z���;0gc�KE���'�m�&��Z,s�,�)Ҩ�K%����1Mk���l���LSkM�~�,���6��vX��-��o(
�Y�	K�p�>i�O�NS�lP>�����'��4�y̝�MM/�mȬ$�mˁ3�n�K�(A���7LV�'�Zc����q�|��k	� [U�˰p��j�	�1/�	�qt/{2��rS������]�|[�!}3N�뗶�6���/�k/�P�a��6�f��@� �?4�x��K�;��g�9�J��B#�z�;�%����j	9fY�r�}Y<�f�l�Ђ+']�]���V7BS/*݌������N�5���Xc�\�0�ӗ���͜���CF{X�:��u�B:Z�LW�-%�NW4w8 $Cb�ԥ�v^�;���h�Պ�G"�V�8rE�Z\�U����}��MF�8����܎��D��~ص�sE���.5A�&zg�����[a����l��5����v�{#nԉp��2|,��B7�LJ>ϡ, �ko�́n��q��scd	���0�2���2	�V�y�5ڊX���V�7L�.�hJe�����:F�b�)#qy���p�(�~O^�q�D�
�u�gC߉�G��u�`��f��n��� @{� ���������r`cx�DBsw,6E�x��i|̅���m��Z?Ĩ�Yt�E���q��?�=\����?-KuW)���I��hG9.�?wS�_Py�K�?ee��:I5\�-Չ���P�^Zڳ4�\F���t9�UH�?|�<b�$�iiz�K��^JM��ǌ�6���\�e�i^��C��Ҥ��7�H��Mc|O����mH�sG�o�9���*�r�o� ����V3c�KK]�3��sm�66��E����RCS)��_diK,�`P����H[}:l3"�Àj�6�l���g��?��jp�ۡ@6�֎��A�`�^��i�&�����酞ڮ�ȱ�2�I"]�}諐ީ����B�gU�-%�єo�e�V�{�ת�J*"i�h�ݐia@�ȐS[���9H�u�v�U�i�D��i[g)�JY�Iw⦁��̇�[��e�pF<#72F��7D�[�X�_۝�
b��j~��4���0U͵E|����3�������|���BHS�(	*�:�K��?�ؖ��Y^Y,K�zU֤�MJ�*[���ԟ�a�T}��8�|spS����>F��O���9w�\�Y��h��5�߽ ��=�c��g�	��SnzpG匢-ee�|�5�����]�C��UA1�|��iSV4�X{'߱߳�XpR�3(���M�Xh1~� ����� ��z5]�sj<kߔR&�HN���:�=n�
i򽆫a-.�P�l�B��^1���M�g��b������V����V��������cfX}�2����7��a����)v$�*�P�������+;X�უV!���k�q]�����`0yl������4��4�����Y�������<��;��ϼ�*�-n��HHFL��?�A�\�pi��x��.cSy2^�`�����R���Y�$��PNf���S��r���TbW�`�@<V�N�=�A�*�zGb�Tٙ����#�X$k�˜b��\��յ���R:�
�XLh:;x�#��BJ����,7�s޸�r Β7��.3�zRb1�>�(1%;��g��r5�_�.�����/˨��9�s2��� �_�A��buL�;q̴�K3҇���ۼy���EZf={�D�}�"> ���C�Q���)٬[
�k�x�i����&e6�	���W%#.R�AڋȢ��5�E~��gٮ5�l�?��k2��6[l�9��G2.�nAvG��L���[���ß	[���>HzD�N�e{bh��}��c�Z���"k�%���"�8�mԶ�L�r*��-�_�5I
�~���衋�\ؐY�҂�i	����PVI�l>�^x�l��r"p�������u�P��W�W9}_2�ʨ�I�0Õ�Ǝ"�:o�{m@���Cw���!�o����S/�un	>S0���}�4�H#�"{qcE%g~t�Z���
��V�8\�gώ�l�:*[���k�%�:��Wn/���Q���I��ŝ��m¶��)��TY[��4L{�5������F(?nPp��X���^��@)C��ה�R���կɷ
�%��%��t�^Tk���K7E�^��z��eTf{Y)y��sа���H����+%������F岏���v֝F+�3����z(�ן��Ɂ�i�W����Xh��XḜ�A�.�bD^��K���ʤ���F���i�{� �L��ه�O|��+2~��2�
PTf���J�˛ڑu�a�^����?�콓����2n\��JL[���&���)DS��{��~	)�q��x;�p�~U���aRGЄ�3+��d�8�d����!7��0�z���72z��Z�Z�*�zE��7�3�=t��6����qU�)�&�I7�nB(d�X�\ifot���O�xXV�8u���ze�U���&��1
ޥ�[I#$�k>�*3������ٳ"�>�sL0f��.?��l�2�]��鿀�v��_��{71�C	˂)P�J�N6��<|���(�����A�0�{��R���q�>��ҁ扤R*��|���9摍m���5F�ڲ�?V��P��}�́�f�g�^��rc|�I�`w��y�Q���ilį���ʈ׉_�b�@�
yХǛ���� �|�2 ms���,�[�����-�������V��@��)��לxtZGo���)*����ۡHh�Xגd
�����G�>�"J��E��]����:-���]��V�SF$�	�X���c��eJl!�C�C�j�0i�:��n��ƈ~A��̈��eu��'��t�P=D.�D������� �-�S{Pj~����hB����� ��ħW���#<�!�8���^��1�Y2~a�C��?=�o�32_� �xb�e¾f��.r�!w�aO�2b=\Mfc���l&�e�x���*�0�`��UH�e�*�E�~�&ʺ����&�8b�(9���>>i@��P�Fn�Ugy�X}��"+��O˴�Kَ"l`W��(N~e4zj)�0$�����M\��m���Dz�"��V&]��r���r��[@���%��k���^�Y89�VO>ǽ�?	��^�<P{��#{�V��fk���$�|sN�����6W|c�>k~�O�����"o�	�A�y�>z�H���d@��
����x�R�#@�AC/��������l��+�%]�I�_#��dkU�	�	�0cN�=߅e1��w
�D�~��%2���$��~D�	��hqf�3�o\�g���7�S&�#5Ɉ&H&�AU��"R�K!Um�;;��mEa��۔O�w������x�Ц����״.�;��d��R������(�Z4P�\��ʱ��̳T#���x�|��3�+Rl@ť7��vd��ŕI��@���s��z��<�P���v�I� R=h�H4��PU�p�s6G�$�`�]p}^��:ٲ	����=S%ӂ�����x����q�ԦNaei%�.�!�U�*�,ҥ���6����z��z���dzS9�G_���~�9�9��F�dwG�B>���Њ3�j'����	��	8�������(0�#�GC��^\��j�dl e+���*�Q-�&t��H	�w�{�攪�</��nҐ>�s����O��Z���d�������?���|�O��I_;-����ؘN3�)�I~�
�Xnod o_�1�d����f5}񂧝!�������rF8+�"������Ҟ�3�p˖|�M��Џ/�J�Vn`CY���>u��1x��,<� ��Ǎ)������㲢F/(�$�>�=%ܦ����;t[�2둤�|��P)e1�jZT�B�ಏ�Z����v䥭��DӚe����W�k�>Z�5k�]I��Ǧ�VSQ]��e����S�
I���6�حX&�N8<�7�����i���b&ϐ_wd�M��6����̘!lj)�s;(yLH&,�/dI��ï�a:�x�86(�[�zx�Ŏ�%4K��y�p[��$ɚ~u��7�+����p�8>�;91,쓿�izU�W-\�T]�{Yl�}��z٘��c�d��.Zu��g����Ӕ%�����?�����]�׏���!��h�]P�{b�+�
��P���k�:�|���7����69��q"�\�V�;_$�r=��ηՓ_`�Ҩ:ʱ8lee2�j�p�M��I�����P�4ǪFqѶ�A�n�*ک�!���q������~�Q�ј�6�؛�G���co��I���]�����v|���Z%'�J�o,�"��?��
 ��GuO @Y��RU8d�[�(�Wh5Z����ުZ�;bQR��z�z��TH�IB�
����l\���Q9�T��[	���z�����o33)��� ��d�2���`�AE �ʵ������q8m����<ݗ��7�)�W��n�����lH��<\�����_����y)��(a����-~��<]	����������X�mA⌙�qAg�/�x�r<�h���y�8�(��U�F��	X��K��l�y�B�pnk�P�e2��*'�ڇ�k�p����˻s�NyS�RU�:jG �Q���p�g=�p���S�;��o��~��MM$�Q(ݺ�ܬ�Z�=%`+σE�>	�}H��h`���
�tm8���;<(����s6�&�D*Mp�&�y�tJ�{�ԋ�N�׮�.uL5��m-*������f3�d6�ad��*�������-�T���"l���m)O/��N��Z\��֞�h����X�X⣽됒'�X�����H���I��M@r�d�����j���&C?`��f����#�/=��M�Y�ۀ���Y������d4��!ZX�Gs�����F�<� �M��?��֔Vm����o\M�Vf���Swכ�X�X^�x����EG�\j�����D�l� �$&���n-_X��,N���g�$�"��v�Gz9���E^Q�i��\4��6����bn͕Pn�����F��	�O��ڧ���7�C����~�k`�4�9�x����Gf��w�^�S]����"Ǥ��P	��U����5�4 :�v��Y��bq�6���4�"�ڲ:S�G_|	��A��<�%=��S�qhd�ͤ�pn�=��?�]Y���I([�NF�}d����m���|Dy�"�s@ ��a"m�.�5֨w^L����n�U�Z�j"���4D>W`g�~ʆ�����YtHbr��T���ӍWx����sȊ��~UL[��Q����q�3,��C--^�O�fx�V��{oG� } 3ih2d!!�x�`SױԪ�ς���p�𡾐-���x>C6�t�fZ�B��<ĉ�V�d9���)�,O�0�����~�wDbͳ��"gz"�&t:B&��$������;8N�a���4F������^��!?�8�6$i�3�W�('F�]���?p��L~HJ�	��-S�,��֙?/�io��'��L*[�:M�"��/�XB�/wV[Q0G={���Rr���%
��7�ܔ͝��Q�T��l<�`������]�VHi���F��Ϯ[G34������\��(z.8��6	T��3�Ed�Q�l�^H��QUSC�g���qŞν��l�M�hh��P������E�RDC���*s������ j�4�s*��Vqc�sz<訂����+�Mۙ)��un��:O;$��ϟ�ߵx$S}W�D9)���ÓZl}I��H����s���Q��g1���/��V��o� P�Vt\��gI�?�S�r�X�U��s0���r>�-16V�/�� O��A
����Fu�7.g��>���R��m��9�PӐ6��$di�W�H�;E/��1�1�dK�p`Ed�]���'����w�ɳzO��Mi/�V5���*VeuT���Y�v��)���[�^��z����~A�̿�:6����i���	1Ȣ��z"ՈZ�g�����<t*pSD&��Ѣŏ�Q�����(Q?��T<=�o�ܵʹ+���޷R�L�U�=FiE�������`�
����~�a`���-Z��%���a$��n�`}�\{�2�v�T;������U�������Z��S��l���9AU�d�=>=Q�Vm�������
��+�:��3���o���^���q[~��g��&�O`�Z�\��o}H%������'�ֺ���[��>�)I*�l�uL�eqg�K�G��)�Q1x&j������y�7�S�o�v��P��g�	D��;��Cvg	X�� ��B�2����>��*�r�[Ѽ赚D��n���0H"r��<дqX̙�
�c������m��+��pUH����p�,SX��>n��n��g��MT�P�/�ص���m읛��m+e��e��p4|�HQS	$���6!�#��헌@~�U۩o�{ �ۃ�����gm�&�����'���D��=K��*��A{�F�ˁ�>3��c�I�wkrG<���L�g�4�<����ܣ�٧�BŢ�]O�X׈F��
Յv�x�~�%zgM3�_�ki����Q��D��{�D�[{�ų�����d�M �@n ��722�Ƣ���tڵ�%�*���R2~˱]�����r������� ��GF`�}���cW�)0�%y6�7Q,[���$��C���@�K�n��U�ϑ�f���G3�r����QfȄଳ�j]�60�;勲�lE��Dn��`j�[#����x4^'J����Ԥ/�^�a9Ƀ�+&8g��!�"2��=J�5�<��"���*[�:%$���viLV��AR�.�,�3GP��� ~�,$�wt;|�g��űb�|���@9Sԅ�kZhJ�$kh��oZQq��;�L�����)����.�{-�%�2�=�s"*3`"����?�6��~�J���������;K�$��*���N�v�5����]3�?Y�6����������ht<�i�Ы�ӚIpuv�/ 5gl	��7�
�1���Q��	Y���l��6;/�C���l�A7p6)mRm��{G+�.� �7���E��~�c	�'Oh�>��
�M ���w��BU��3{���2\�e��0�Ɲh�X�LK=e��X랏�v�
�d���_�n�Q;C*�&�5eU���Ty�~s[��^ u	�p#��P���7S�����f=�BB��῭]��C&9գ�w/�
qH��GJ�ufж��ߕV�*^9oo�0SP˗|2|M�����h�6D�Sd���B�����l1��q�RKN��[�\�B!�`���2�M�m�{� �Ï�����2M�m Oل$��Z��XN�tO�n�e�7�Ju
2P�-����x�M2�O6� f[����O?��Uo?N��a"��8�MOp�տ��[��F�˙T�@7�=�:)�ň��
�b"ƨ�n�I�<Xg�^t��Z����?L6a���f�,"��5�K��9�ҏ����n���7.FU�b�o(_��SsNB���4�<W�@���p���w�"eJ�]�7h�G��Y�7�Ѥ��/L�62
�W�Ks�O� 1���������M�wy�:�)u�,���UɝҹC&'���<�%�_��'Dk�svN�ǐϤK[:�:�-�baN=IwL�:}4��B�C�B�b���}\����*]f�1>cN�Bc�-�񬶹�ÀQ:��ֹ�|�%\�0&�ゲ��K2b�Q�`V0D�g���R�FT�r��<����֊�\��ƋJq'�g�F&Tx�]&������Ɔr`&
��x��x��i�7��_E�E�U�+yT�D�یu�iE����0�#�	��.�M�#�B�d*�r����tæ�_�u�������g�P��������>�>YF�
��' Z�ƺ��ݡ��0z0�s��zo��*X]t8Vx��v]g"�� m�Zę�w0���??5N�q��-)=�J���r�*D��4A���Z�8&4 ����F`P��J?����s)+��j�*0�.����w�'����+՝ptT
)��80���u���2_���*���\���L�W�"ڎTA+J=0]L��<Q}���) �%��:��U���H�3g��@C0�o~����z��g�"Vř���f.�|�[K(�Iɕ�r�۸rqu���5T,��L��JF]���Qn��} ��4����U����P�]����j�.�ױ�°7{�6��	bO����诠'�z�40Y��_�V1���-��?S�$�΂�!�^���j�{G����M�5� ����Y��x�����V�mǠV�3Me�:��A�l�����F�b����o�@+����S�
�4 ���#X������rW��l?j����@�Y|C�2�tٓ�e>�3G;���콑z�qkNq'��u�N�_�[������#
(XL�H2pM�`~ �ǓT4�m��Ἇu��_;�L�_���5�[ 4�gO&K���^S�x�EˢW�T�	;�ݟ��	���[/���F�Cx�8�6$��W��C��r�2}Q@�֏���sID���6h�/(8�c"ׇ���bvc���(�Y�v������=Fx9���5��v�(5l��9[�(/�r� d����K�Y��+P':�Q�vƉ9�%5�[8�{Y�ӌ��+�N����M�س��ۥ���Z�����*��_K�eh@��$���E�p��ױ�1��O�B��AG�3/��G5���6��t�%c2�ׁ��Y����X�rnZ���6����7]��,��:Ĩ�D���fT녾��4�-Kژ��_1vdt��t�4�}�B7����Bi�Tv�R9vK�E��{��C�@�
�b�W(��Ql��*�� ?^:�{j#�3�c>�u�P(�tEhm�^��J��x)5���)5^���A7����$h7��k�K�|	?xن4�p_���8�e��d�?`h�}9��fI_�*+h�����ߔ(�z�ًw:��Ey���-m�+ż��^y9s2A�S��Y�zW�}�t��ƗT���b�~He��� z`1���Y��9�k�	Rm�kw��pfg����X��L^�%�v�T�i�H`VR�����2��2�*iq�ks��^MX�8|k8����J�P��kk�G0E9�|gP%������LU���vA{'����O�����2����q��+\��Y2g��C)`̅������)p�/4r��BzG�$�>o�v��*n��>��f�]q^;'��^jbO7�?�(�'���[X��d��)����̱Nc�m� Ȗ	N��[2o%3U*f�Ԥi�Y��g�.7��O���H�+��	[(�U���㛎U���/�f(KΨ��W�":���px��N�c~~��L��CHٓMvZ�^���������T���Z��{[\��2ҟ��%l�o���źP-�̥�r
��@���纑����<�����(���61Q38$��I�v6w��ܪ<����iq�N�I�ogF��I��V5;=\lI]��f1�G�XY@̃8c^%���`�=	���u0Z�&�������MĹ�Pvd�1���G��N���:�s�\|��h��ă|��&,��_��Hģ$C��te?Dj����G�~���y��KON�#@�J�<��.����Q�`�_� �Q�C_�t�kf3��݂�5]e\��L����a�������dy�y�zR]�ͦ����%�6/#���|�D)C�X!�d�
@{ײJ�YR�w�x��
�`3ܴ�lZ�G��M���q�k�A|�,�LDhؼՈz6�N�K��P����sQ�|���~N�&��zX|���}���hh�@�{F�Q��o�s�@���N
�$#�_o�˕ f�l05P��h~�ʚV9�|U��i�cG)��l�O'��T`7��� (W@��ТF���b���T��� ��z��t "�������P����3텬���k�d<��c�#b5v B���57�P�麘�`��7�:����aY+�T��	!�ʨ,!t�x�5û/s���Q� O/K�1�!�?g�~"��Z��qa:׌X�!�pjP6��Kr�ΥUW��>������S�.ѭ��C&KM���6���y��"��V;�T���`_i�����ɖP���;O����lWԬ�]'	�v(7U�L-���gP�b,���V܄�pw�����2H���|ޖ.�����+�I�_�����`~~�#/�50�?���X���J$M]Ngd�q�0��Ӱ �.����O�G���ӛ<�^9=��t�`�;�t�_�C~�҇Ь���B N��'O�z�;��L�)�	E/�	HV��Y�L��1�)⛦��'Z��~cx��*�>׵M�Jyx��?�
����7��P<��c�j���_I5��ZR��k���W��:�{���������|;�,7�����T{��6ǵ ��lB]��I�
25N�3H�(�At�DcY�vI��ߏ��s��U\�(À9���i���h_2�f�'ǿP$�UG1��Ca_i��v@.�5F g�k���tnaħ�b��m%��_�"UƖj�����
�7���\�.�l`c=*;�Q\��9T��������,�4���)����a:�rKj��R�������/3t_�N�i�d����ojJ�O=0EB�)U�Z�������9>բLSб�]]G�A����� M��IЊV^n���$Z��'-?�:���ʖ��A����Q �8��H�˰~��W<�6hk�W3iݪ,����h=�C<O�����P8�7.�9
��-+6�k��h�p&yf�V��]����(��C����K@ �jp���tk�����t���p���"*�Y�ǳ�9��O���PXT|��\�Dj���L��S	
��hez(��S=Qɶم6������W���X�|Y�����󩝪`xO�@�A��$��B�CM�� *e��%��NlѪ&д6K=Sk��/՘��	}���Ó�ֱ����Ĩ���.3_MT�#�?]ĉ�m�s!�+�-�O���?�h/kZ�_�(7]��_ �2�5�k�:��JW۫
��t�R�m�`m� �3P����1N�\����Oع@Qn1��(�^j��!ZH*��FHq�T�yZ6�hK��Oc�X����x	�����%��ԑ� G�X� q�{ve�$�4J��y�����a���K�IsI����{G�Ym��zv&����o၈:v_�h�\#�-k�Q�!����b��� ��j��V�i��M�>?D�*��u�*5����]�ܜHI���T���`jҧx��9�W�&FoH���u��J�s�BF�^�� 8e���p�sO\ǘm���9)��&���c
l�NҞ�.�����Z9�h�X0 ���3kTlDf��}E�e�irq9*Ҏ�kˉ��fc��v�(�M0�_��*N~�s�g��p���$.M p>�Z�x�,5B];�'��yH_�Ҍ�m���,�*�uu]�l� 0;��Ou�Y�-��;b)�Q5�dN��V��z�ʤ�x{p��f__n�g��E� a�r�zo���`_��lC9\֗���ֲl.>y��@�>�n�b��;s��"����u�Lb�ݗe�K��#��^��DL���N��P~r�����[�Z5�ʄ�4*g�����^]V�b8��c�ɡ饠��������-��_kt��G�>�����~
��Dm�i�
�~ȅ�B���#��������mу'�	B�`�U��v��m�N�p��h?7NT�ya��([ߍ<7(q�M-b�"0���N*_�v|�ʚ��P�O�F1�j�ϸ��j5��������k��Sm�g��E��K΀i��M	u`H�J7=;
�kؗ*D��|�Ue�R��a0[��8U-��"�v��7���D�1!^u�@_]��1S������\n+?x�h��w����?sd��[:��m��D�������]}ɺ�x�I&���������`C�
�K+�$Vo����Ț�HTz�q=�q�J���О�,���4�K�'�h�̐��=���Ya�M�B,ү�f���}����޴w�:�A8�Ũ�yz�1v�SZ3�$��i�y�k_�����o��aL%q��@⇁��������F(䍰�z���7�Ӿ��@���j��Y
��(+4�ش�c�N���Z(���Av�et-�A��?z�oE%[mBta|Q�&l+�åH�r�������(��úJg���X�7/�ٟ�S�H9u�o�w!G79����>d��~��~s�����h�F0�x���Ã��G��i��|���#��-2����Q���A ���/?���~��0>���:�	�����@��Z{����{
1�~��z�p
	{8,�//�M�Ƴ�D,��6�k�*댥�t���1|pЗ3�cBS��n�����O�*�A�,YZ���L����D�k'��+�����A�J�O��Ʊņ�Y�-��agƣ�D�HH�Y>�����p�*1%d�06%���Ę'��S;�È��4�+�x���3_��E
V�6������-����l8�/X���qo6^A5IH�zY�}��J#X��i�ֲ�-�!�QBgoD+��1rPP����#��s:$5�2�a�Wd�;��)o�1��(^��haH�@���$7�~u�����J�k��D�-:��i+�(>�;���`D��у9�������g�-V������2*˘�ZY�4�0#&d����w]�e��R���,y3}>W����ײkX�ڪ�b�ś�q�zz�L�3����#�x?��J� ��'�c�N��f�����:٥wK���@�zqE��s�z�U��5���o��KBR�Rrj�L`���4�����a&P�# ������K�8c��ģw�����halԉ.G�¹�l�W�D8h����ޅ���j�K��@GXk,����S��I�����smK���ю�%��n�c�u|�o%ܙ��(��&
�p�:�3޲�~C��RB'uk�Kn�6���U�L$�N�O� W<!�[2�K
���{mU2��Ce�(�y�U1��Z˦�8��aeFK'p���EE���RL��6���z�I��c~*�a�.��:i�p1�/<��#h_�
S���s�f�u<��-p�GE����Du�������H�I����O�|	r_&�Ws� V����7�4R�����$��>Z� �����J���z!��~WZ�A�L������! 膅{{)��Ώ�� �
���:�쓤g�TM%3��C��)�l��y���i�ϝ�df{ey��%S���[zn�eY9�yv9 Nq�?)�D��^�&�2+Iw�!�/_��H AH˜qOM mQ5�9U�JAOh�%��C�ёA!W����{�5_K#�<G!����T�R�Ѵ8^�-�8Xm���K�����zO�r�������۱��pB���c������/f�v[!l�J�����9�_'G�BmeZ,���.�UUU;�ca�By-oR,9�X
����Ҫ����-��;L��E����2�c�w�,B���@�M� �����X����y�l�5?���K9����^��ǎ�C�����6�~��G�]��3��U��j����� 4��1��#r�)\z�%�	el���6��`^y�`?f�!jܾ�A�01%��q��8C��`��M�������v�w/��kN&v\u.q>��, i4��/Sĉ��z��d��ѯ�@�u�P��c�I}�B[���ìXvV ���c�3���X�O v�;'>ح����$��<��ȧ�����'~u�lb��#Y����������J���9��4�u�4��5��<��;5����G7�H$� 2ű7U����}�FA���<�()U)nuf/�����7�*^g�U؜)���u�a�+7���[�ʞ3=A+;]� >F�����cq�n��� `���h�>�{Ʋ�!�t��
��_�PLC�������|�M�����wv�FM!@�{�n�����\]���t.�@�>Jy���>�2^�r��-�|�(�.���J#���ﳐ���U�<ګҙ3�~�YG���Yb�5,tg�y�f7~=-��'�=�Sp;�Bs�R�bK�+��o�s��G��AǉA�ͅvZ;L>��Z�$�/�ٟ���J$'���4Mzu��i�� dد�>��Q�r&\P�kiO¿�g����b�޻D��K��/=�띪.�@�����q3Oc�b��x�36X1tx�.�G�%�yu���K�u
��K뾪�O���h�S�=+:�۠���EB�,PO*IA%��槩*knY��A�:��'�&Y�!n�	m��y�|u&���&wڣ<�Vh�r���ԝg�=c�XͮA��,��އ�e"-�!���33@ڭF�Z���/e=h	4��dD��2ǈ�����L�	H�>՚�}��'X�~;�n�*qâ�t-��x��mƾRD)�L��ΛoR��a�mi�t��z�1�����(���)���7�6e�
ۋ��8Ͽ��h逭׀�$�ܙq`�蒪�3+�~$�. ���jB��:<�=�$&T�/���a�9�R
s�p|��S}�k�cK���|�)I� et����n�䖙7�ٷ��*t��+�eX(Eop�0��'9f,��O%��28�b�"$p;�{����0;�"�(��^.G]��h�� ��W�	#P£�X:��.�C"�<1o#��.	�8��6�����F�o�8�s?tw:�F|Y�氾֖�@�FFm�C��p��n�k�7`�`��B�$�)M��@�Fi�+Ӕ�{�3�Ȱ�X�{@�������aύ&X{�F�Ju��%�H���ӽ&�"�5+z%B�Z��!�]
Vowњ״��V�A��h&�;U��������w�<(�h�z0��{N��|Y�N�/�f�~��D������K��� �X�5�	U[�42��o�X�䱺x���xG�vg^��CQEm6�^^R���/��np�>���#��i,]S����eLe^N�#�?3@�7��d&]� �j�*5��)��e@{���{�Kl�QP��J�8u�`�?��U�v�:mo���~�J�˵�O�C��S��:�;��5�Ŝn���:'?b �2&�M	S���FW�P��$���N9�Z�
�̐�Ⱥw^�P�z�X%C0���<�E�j�$��z��f[�HN#0q���fR���'���n�Y
4�e��� &K�e���Q�����%K���+_ȚQNWQe�l�� ��Tn �D�Kf�2&e�e��n*{����-a[���jh���=���Ӹ��B��SZ����O\1hi|�^E��<|�f�6�^�Zِ�b?�~Ȑ��H��:F��_��f�p��J?3ѯ8���l(�L�*F7ۭ�'L�vn�/
����Tfm��rO��n�*�������Vn\$c]�쀓j0�e	�b�"�=K��=����J�5o��+�|h~z
B�+�Q�4�	���9c&���!v�r�:���A�9�Z;��@�d��#������s�-_�z�"j=iBB�^�����R�v������>Y3#�թ+��]�]8fkZ������q�d���{]�V:�7q������ ���~%u���jDV����/�#���=����M.���@��OH0s�Xɹ�`�> ���	��#�b��|���F��֌&�?6,y���a`���=����/�N�j��1�@��1
;��F~6�0;�*5�%��Dh��p(07���FNi��3SQ���?^y��z��{Hk�{~��俩Aܵ �d^q���<�9�2C<�^/��%�������2�F�5Bة��i�=��wH	���O�[����3=B�G�=K�&�FK+���G���<��S)B�Nk��1lE@�3=@��|�R����η�t�6��˂`L
��7�,ֻ��#-j^���5���?��/{9Y�&�|/)3n� U���4 ����i�:�KN0�(�'$NC�;�% @.ҷ�魿,���c(��r��ҁ�D#꿞�,u2�~J�M�K�/���ݭ��0�V�"���D�+�ZWG�8���zq�D?��v��u@��U��(0� ^�i�=�&]��ԔU�f4*OTF3O=��u�-�d�iZ�jOR������f=�<�x�+#��=�p���v=�f,�`���䏀_^�Z�.�� ̌�I~��Kk� BO��U9��R�5\�.�x�W5N��=boM�|�� (u$��s��2Rec;min���~���f�����XK+[�I�n�{�eB��>��hTt��;����������c���-ңP,Ϳ�.=r`q�A*�Dcl8�'�ԫg1)�䍗娀 ��ڜ/�n�����ٛLjx��w�(��!G���e�덳���i�V�H|Yd�_Fל����M�
��d��1��g���g1�ϡ��(�Ox�����;�� ��BG?��&�A��/h~-,����v�/f���KR�\��H��rFc��ۦ�i��B>Z�u�{ˈڥσ�ہ��@�2:˴߁e�y�`��y��J�!�Y~�`�U1�Ӿn���B��q�Zc�>�^�� :��
�<�w�� X�{:p�q��1�L�ѡ� v8�Jm(���9�9��Uq�>Ӎ�G��z��W���]�wº�_͇�6�����R�R�w�3hY���r& ����������3wN��q����B$mɨ�F����Ʈ�5�!atz�gƯ��QN��@"W��q��`�ȣĝk!�҈�ް�ΒP�������BQ�A�k��)��%:���������<\).]����� [��>�݂�	��H:���n��p1�K��m�GW�/�W'�*�\���/I����Pm{��u����G@͞�E��ݪ즯��o{�|S�W5yq�j�v��ܝI�6%�ՠ�[0l��8y����Ѐ o���*[�H�]� �D��S{�$M1-58���Cl������Z5�R?e�k�_\�z�_��;�M�#��a�򭐢����0���<�P��G��&��NP��gԃ`�G1�c{�D�n�M~Ao�u�v�4��V�F�$<�%���;�u��n�:�+�H�M�Ye�<����©I�����_���g�91�k���E�p��W=Qw�螚��i3T-!��
A��-��i`�I3����hy;9���ɟ��¹���讨��7�E���}��E�?�������4PYx�3��XSx�L����|��$I�8�	P~6��(٢P;�e,��ϩ�M��R���1�jr�c�,ɠM��Tb.`qș��0�67Oa���g�x���`��KZް»��B��YC�)[�Ŋ52i��T�XO@�3����@¾s��wǊ�M����o՘��w�m{�(l���9�U�0��NU��W�w���͛w0���.�Q���c_ڔ'��FUR��Tx"X�uC��g��{�T� ���JFRS�5ڸ�GLI������v�Y���uF��N6���1PX��gy�a�S���z�v��|���K/�Z> J����I�S�T%:�E��,"��@sۛ)��G#K' �7߽"���HC���c�yŬ)^�*T�� �ϭQ�z�e�RPP�<g�7���.ұ3��_搴˺Z;��|%� �Bu��-��ڤj�؊�� j=�lk`Z*ʠ�zԾ'�gk^Ӹ|D�� xF{{�S�6Kƶ>߶ږÜ�}#�'��<�_��A�O?\���dn��kFY��Z���D�s�,�ؕ�%8
]�Дm�T*���
��8e��.�����@� tDb�΄龤\B�u��܏�Ը�r�:�un��KP�\���pu�M�Ɖg|��;�h��P�s#�W'4��]g�� 1#�:�:}P�, UI�%1��ff��s1q1b�7���I����5XU��@�.�ᳪ�Л�5���͚�UK�R��R�oꍯ�f��5/�,y��ҿ7��č6�v�#xa�r��N�H�] br��z4ݕ��!�\��
a���p]a4r�].t��J�#��8��M?��p�` <��]���{�^�^A��?ě=h�D)y52�j_�Ӵ�/��I��Ě��Yb�/)Į��t�k��dמr�WloV�`C��*4u�Sey�J.s��RČmL#_��O�}��� ��`P)l��9Vr��G��<�g���6��>7���i�,�m�!'���7))�퓯!�]cUX�i�'1�z}N#Y��٤�x���O1�8�j�s(�6ұV���B��r��$&�2��F3�즙�,���>'��/:���o1�I�k	�جD�;��۾d�sA��<[8�A��y���>7��>��?�
��/ w�ρiQR�o ����ܴ��É7��<����y��X���Bw�Ex�oE����A#u!�e2��������w�Y��O��Z��"c{_�a�C����6��k�S�p��赕�bV��.�e����j막��/J�<�t,�T>�kP�%��@����C����p�.��;ۼbƘR��P�6�|VY3?��(��G87��<6v0�M0 !qUe�0�62�ɭ�Z���G���[�2)_}+�?*?h1@eo(����M�(k��7(�y�m��6�OH�t�3PfK�Ĉ��PZrM�����j$A���]C$��sx�֋�dL�ȕ{�d�R��U�\�ac|+�����;l�t{�Q���U��OΥ�/�S7~�0����R�l ./��V�8�����On����w�P1���;m��m��1�E�˅:���.����ܩs�;:��k��!?��}z�E�]\�'���qM`A�w�N�Eڌ��Q�nB\8�-l=8S�$Z%7�.�ʆ����7+GS���l�qadެ$�k������2<�[�e���n����W�w��ql:�"*R�!��D����ZyK��k���yɾ����:'���I�?���f8��-�F��w�p.:xTg��(�����+u�����=s���t�M�^��Ns� *#���9��R�6�(���v���߅S|̛S=�}e:aQ)���/zq�ήl3ϵ8v���iO��}Z4�t�rĺ��O�8�"��
�f^���]��f� B>�<<��b�Va��Fk� 0�J}�FVd$��"m�f������'�*�4��� �����{�A�����!�!n�9&~5mS�C�Gg��*�>����Ha��:�*4Kٴag�P��?jkT�Sͦ;�vꦅ�{�c�Z�c�Xܬ�Jz��g7W�G�h��SG4���@����������\UbM�4&��N` ��u�lBD@�D��ܝ�RW�7+�ec~�ꫜlP��f��_\�HA$g��w��񗙦�ö�e�)d�-�[��dN�~�Cߍ|vб�㭪�0Fh������R�A��a=`ߍ.��A����Z�	�7AX�q���l#Ǉ�TѸ���,�����}���[H�.�ۏ�֙�yQ�PA��t�Y�+�!0O��3�?�-���;�p9<b�=/�.��q�ΑN6�+�vzA�P5zf,ӴR���é�훗�=�J�̷0�0�ЊOqך��Ȋl�ղ[�Y�5QX$�_�k�8�VLW���� &�U����v*�� x; J�0���`�r�&�vX�w���i"�T��>d7=�og4�Rd�ϟ�>N����B3�*��e�?q/���4O���<#�E[u�cѪ?�u N�b��ՔC7ubA1 P�h T�3��r���@�ބ�2pe�jH�����bM��D�u*��q%�b�wd�)^���Nhq��:���W?jv/m���\�$Fq�9��R�>��b�նܞևv�hT�$���ӟŏzO�S�+��~�s}�2~@�q�k��DX�Czm�%�gUK7z?�؆n�L��2�[���s���q!������:��f�i,���,�I5/X���F��,�ˀ"*F�qq��R�\�I�LӀU�$�YE}�T1[�l���033�j����<��0ba�}Ǟ����ZVu��d��Ze�V�H��A��þ��#�8�]nf��&G	�`7!��V9�g��`v����� �|[ۉ�bp��ym_QA�1:���i�%�C��h�b���vC2/KM{7[��ml�o-80@ɧ�����{|݂!H3$�FIމ/���5��[��]Ω9���>��1�(�YH�!����c̺��=�[����w`#P��/aJ�ѵ�������Ǽg��Ȭ>h�7�B^�u�"��|�y��T��>��؜ ��ԉ�VXR���S���=�c�@ hN�Em���MV6K`�t��s�G�Ɏ�D`�F�b���S�;aG5W���Zy(����gX�7?MN8[I'Р/A�v��b���5���Z.�A�}=%���f�1���4]���l��N��Ue*����vH��V<��uL��t���0��=�G��*븅�}��>�84Wvo�g�;�6hP��.8c7N����'-3�_���Fe�C)��a�m)ԷH��Q�Q�G�df b����t�Z�P��������������q���F^�I}��n�a����q��}��3+o�s�	,�Q���,����7������<�'1cw "8��x��aZ�� �`ET��1P����?�;�Qv�"�cP��Q��.�N�j��]xk6E�덢3��~��_ѩ�a�O8����6��5�4�p��y��>W������u/����r�	
���w��NM�6��g`1&7T̯\^p�.���r-�^�Q�S�o�2U��M^��1.o`.	�C�<u0y7l|/��ӡ�q��u8|��^]��-�voG�Z��$�S7�դ�t�O=�-N�A��7�s�&��� �솷���[sf�gI�د����g9���
N�(�����_+����'�I<Q�a�{Y���_��i�X��|�3�����x�["5l:�݋Ke6�+R�n��<�,'��o���T���(�kutjFǧ�pt��kk���$�"nf���t���ٽG�MY�d)oRt�C]�	�VsZ0��o�o��^��<�9V�a��s�� �1 �}e��pPj%�-��w!�����YMJ����K'��a�C ����jB2bJ�d�F����ь�9?]��YZ�ؗ�3��+`\bg`{��(�u34eؿbM���*[Axw�B�%-�rG+ ��uTI	g�x��[U�~_'g�k%I�	S�y_�"H��D�$���]G�r\����������g�D�J�Ȼ��Vm7�a,�hHo[2�c�C,�܆�iqm8��k�0Vu"�\Z�c�zI]{A����o�\����M�~�K�uq��sa�ށ/Ɍ��V`X�����r*9uT���Γ��wɞx�Oda������)	Y8�w����R/�Z��q?���OuB����ВN�ұ��W�2/�.������_\F���� ��)%ݱ��(�@7��tI� ���TW�Pb�C��� lx��;��Wrg"g*!�
h?�7h�<�W���)L�o%p�X��R*����P��)nIK�*�����M!C_�r7����p��!]@跽�k�X�K٫��MY�M��/��1Aȗ�÷�9^˹�T����Ƚ1���F)���Z]�z�]�|���q��A�,UO����>dc������[ ��
r��x谌0��SA§�yM��kـ��m��:�w4�]9'�l�4/�����ȶ�ŷ���Y�u���*u��a���U���R��?���"����1�z�ftH��� �!�Tj`�/�;E�M�P��Yyrg�4��חM��F�Ŝd��X�E��%���Y4_ M��81��a������aA0�X�)���>���ު7�z���F���}�(�f��0,�[
jZgM��������̧���S|�l�[I:�k�q&�x�-��dׯF4'�M$j�	~e��z��ح?�cY+~���0�B6��m�9�B���W3����[	��gK��:���s����g  �{��\��%	kD��.�[�c#�d,��l_�G�O�Wf>��
��+����䔍��z��n��7�f$�劮,�L����6�:��:�P"����0'�˔ux��"6�0�E�]��PM���t�9�oZ>�@��g��_"sM��D6(�G���ឿ�E�J��墌}P�۷��j��W��a�(�YǤL��}���M��ilw��)�e�h�
p�1U_\��Rn:U��Z+����[�%i���5�u!Y�~��7�PNݧ�&�f��R���W���	�1);�֛�����µ�*��Y�W~Jw4�ϊ	��K�	��dMq<�Yև :G����bg�kBY�wx��PYP�RZ^�=�o�(�^�]�����Cw�O����=I}��0m~&��}��R����e;�9�T�<\�E]hp�͙��Ы�8�t��*D��Wf�˄����f]
Ua�*Yp*D�]��y�﨡��8��s��Mo�]�� ���팶�^��b�n	�o��j«x���C�llr1w���Y~(��w�#��3�7x��D���BV�p�e��P���_ѩJ�����F��6�a����й�)uq�C�(���>�boJ"������ˀ��|��L�a�LVtyC�P
oD�T:�dʹZ5���8\ðn���o?J��3ݍ�߁鮼^+��Z/	����ؠp���5�'l=��H��9�����ZcWՈH��T�4ᶘ���q�v� 䮘:Ҹ|�r�Sͱ����֝��{��d5��0�ks�חs�^�g����V�*']�CP��[�����\鹱�8�	ww4S5����u�Oe��#]D���䶌lx��wF�"m�zkC˭Y'�\�'0&��fske��!O���������P���D(R93V(S�I*?��.���|��<r�Hz?H(!t�Ja���`� �S��Je<�����oo��-�}��+����S�L���4��1���;�΃:�1����i*y��0R|�A5��-�X&��i��;��o����3��vǃ��Ш���L�V�U�ߪ�g&kV׏e\��~�����&�K�Q�X͌��/L��N,�?��_�� ��C�Bs���Y�c�<�ԝGlJ�ߤ!�����q���V�j�5v�2��k�7ښ����	�&�t�	ڄ��5퐚um�1��({9f7�>�S\�Q����W>&m���}E�S��9mC�A�T|�8a�����Ry*�.P�}�퐠�L�,W��Hvq�+0�����H����&��jz[��=��\�Ο��CӒ��!Rd�eO5��4n�S��ѡ���uX���65M�0X��60�W�>�ȅ��U��`�Xy���і"֝�t���Ҏ�q]���o�ؠȀ)T&��0�4v^�"�4�A���>7e�tI�2�c �����r��X�BХ�Q�mN�P��Y����9O��l1,06�1���[�:v������W*����H��R$ѡ��`P�A�6_"���=d�� ��2ᘠ�JG�":x!��S��c82����%T��nH��lf�o]+��h�I�칭�6w���N^O��P&ek��e{�8}$NA�6�`����|R�!փ��$�$#?�3������r�G�3oJ�Mm����C熨�U� 6y���d�3ԲV!F�6ƁxP��9�'���A�մ[��T�6P�ʅ�1�S8Hz���^�&�ͬ�uJԟ@zӆ(�l<���H�����.�!�\�h%��6���c���ƴ_�h����7���<g" i2������:썍��6�
�F"�k�~�����'�8��~��np�Y�ev��J��|��_����4
�#�w9}��;��B6H$h�S�l\5�����C%�L��M���5U��CE���M ����h�Q���i�i�x-vb����#�Z����Y��E�\��l~ߖ��jF���T���Ƀg~q
}G��L(��%�m�U�D�]$���P�������������CgĎ����#B��{@M(A�X�4k���9�A"����v_+��'u>�8�vW�����}�ᴡ�.�R�(���������3M�,7��6~�}�P*����[�0)�j�%y�cyQ�4�M�2�$�kX􋂛(R��nW��z�F8�X�I��^�-�c�YW���D��d����m��@�)�E~5"@K�ڮt[��Y�Ԑe��Ih$pB�k�<�5��x�u"ٜ��4�2qޝi�7,�v�U��VH��<�c{�Cᢙ@Q��
���7ӛ|[���@W4��3�b��7mݦ��Y��?.X�s?x����˯&�!�=���|�[��?���n�Z�J��>DU��Z�^#�g֫^�W"������E\gG\?���"�X�@@����=�A1
/�ל�U������v�;�q��V) |�^���~�NuX�ܞ�n���lF�3�C�Kz�<��g�9߇U�j�.�PSc䃇m:���]�m�83#�*Ǚ!N��zt@�?���7���'-}L�܋���5#\�L�H��,&�jη�#��3`���@I�D�'��j�O*�U<�����1�Yag�cdη(Vws%h�n/�L+�<��[�ޢv��Ə������+�M��(��$�S���ܑQ]2D���i��e�|$�-/���M!f˷Z7�����T����Ƽ��S]�4ם$�~�b�l��Q�)�'��)v)0�;��[z�v��<I
�	W��b��JC7�����c�2���[�V�-(`P"�q��I�k����ۑЪ2�S���W����]� NSW\�jhh�Q������-�Ń�Ą'��A<��0ߏ#��,2=��2Ct��W�̦B��j�=H�V������knLZ�(B��PI�1��,r�j�-���ҵ�	�0)mkO�Y�Ƿ�6��^>-��5;6���2�}(%�l(��r���O�i�*�B�V/����\�)}�P}�}'�K(e�ݭ6��K�IZ9�!�*%p�Į��R����~�[�e��x��ծ����!Ba��M���@�{}�d3k��g%篫�m��ruʨw�H��a��B����)?q��!0��w� �O�0��Ps�����F���⥳����3�.��>w�8����C�jN��6O�~䅬��j�[�FS�u���U6�@:hÙ���v�iݡ����H��\?J���nU!�?&�
)���:����<�����@�}1����+Rd������O���KQM������LL�X���~�!p�<Pp>.�9����lo�3����t\�~_�����%��*#{a���1o*�v	I�R���f��:�GG���N��[��ϗFn��)'G�MD,_Nk`_~:Gu�����WQ��ç�#!,���I�qu�/�o�yVAV/�*E���x�GF�/�_�T���*�ҏm�B�?�SO����T�������&&�2j	?�x�$K3�n���Z�=��<X�O������	��+�����l~ia�_��m[N�����t%�L���k�+�R�ɔ��N<c�{��|V����������[u�s�n�J!��4�����LW<<���7u��f�~]�.=h�O;5�,Q�
%NL�'�Euq~�е|L,��"؇��7��Д�F�Q셕�ֹgN����39�b���{Bv��D:���(7�;XA�;R�	�Zg�06}W��h&q�}*����yt+Չu�l�"ؕ�ƻ��v�6�^��P�8O ~{o-���%��2��[ �8� b��VK5¨QXE��ԓ��)Fέ'ey�]1����	q�����qܝ���D֊�/��r'���V�;$'m�P�������7"��5�ճzt�c&�]�ڀ�!��kT7|��}���Ƭ����k���N]Dsg3�j�/�ybr�.����o<�	�W4��o|N����G�^e�[|�Ǒ_eZ�}*u�<��j�{?��R����M�x�A����*p���.7ĝ��ٚkI�݀���oҮ`�B�A�QI���M<�k��G�����Ԕ$�Rɺ���g͋ﳄ����6�!�^�8�6	PE��w�D (���-��e0!Y�O�ݹ0բ~��+�)�g��P��#�i�jX� a�Y�=(r4 ݚd.��R�? Y@1�7�)i��o����RB�8�G��-?'��#5M�uL#��%��}��I�aIL�L�OR��,��%�"���uj^�N�eUD�S߽�#����-7H���%�y�j	&�(=�k�>����w�U��D*3:��V5�yG����-�'�s�}2~�_U� ��Z��;��^A�z���|�`H�~�;ܿͭjxf�S1���m絳�@�r�5�7�^�|5�M-1L��g:a��m����nA���[j�'s z�*Pa�8�,Z�N�A��"~���S*n���3a�����1�fMGqu����
`e)��S��'�R����d ��l ���v߈U:��LmП�7�b��V!�90�TCC�|W������j�8����A��m����z�P�⎃c�F?�N8�p���F�sj��T�����ɫ�:8Ҫ5ʶ�@&D����K���ԍ������l�8Q���z) �f�~�$V�Z�XE#L|s6��Ab�
�3���_�_���t�v,
���4v,�0�®��ޑ��7�J���e��P�( �3 `/m������\�lZ'q*ZC��L=׀,a]�C����i��4��{CZ�+���AO����y�,���fh"��y��5��(���+����������SzXfaU��k�),���X�q�{#���aa��9WQc�t���~�<;�ROuRv'G��]�ŷR���$��6b��E�KU'Z�&8%;�'ga��Xע��z=�^��y�uD�|�_�Hd���M�@����<h���̈́�\��b��7u+�ß=5�r�֑������sg����4ie��I
T���؞�h����,h�^���m��[n%ts�i��5}	˵�ia�sd�܈�O�Of/�S��=�<��Npu��b=_��ٜ2��|�μ�-[�?u��k�\�ϔ�OV���)o�����B���O q6aQy��w��y����xZ�-⣶�U�8B�	�:t&D���Ǡ�Ɍ�u@�����3�ڑ����/�3�=�8���b'�'!�7�Q�p�Æ�YH�	<nq��I+���qv]
B"욋�qP��f�&��S�ujxƍ�*��}���,���L(?H�j�B�l���ǥz�EAI�&��^$_���c��ٱ�/���h�߁�$Ov���"<�|����E�\�8�-DAW�A�3�S���k�=��뺸� �W�u�7��a�=L��}�o9)�^4�j��0�����;�sl��(e<�E�R�����e�%[z�-���
���-:�%N(�Fٙ�+�#<
@e6*?��pR2)('���0s��v��V`�&�+�Z� b��-��n�K�rZ%_X�#���,��Pњ�kZ\,I[�H'?�x:�K2����s�.g���6�o6�C�����k�鿣fݗ��_LҢ!M���u�ܫ��������O����>���H1���\�K����s�٬q6�/�~r)�0��=�͢����3�9�#���ja���t��)��v�������XQ�~%B�-O8�MT�O�=�}�2�҂i`q�|-�䌼��:�"���^,.&q��ݔiW�f>�иz��sn���Ŕh1c�pʛAә��	���3�c�9:Eǭ����� i4`���]���奢"i��pT'mm6�iY���Y�m�ּ��d�t�L����F��n�(K��W�,i����z��#yliT�A^N:��#�|&���֡	G+����O���Y��U;W�2#9*T�q'�$Z
QpM�c�k��S��r'YN	T2��8m�����elѝ�g7��*b�l$VB-"�PL޾ ��YXԥ�x��%�'�Ѓܿ�E���i���i���r�?$�'�q�x�+#X$'�z�ނ���UZ$�9��D���w�����څ���K���IN[�Жz�Zm�F%\���e���@��Ag�F���bz�֗���dj$�h�+Hq����u��Z��Ur�s@b��]��p��xƮQb���*�zN��c��:��`��5�g����0#[���z��N�|��x\9�R��L��Ukg58��|�U$�Tk�j�Ԇ��4�z�L��Rc��렢��������qپ�ؓI*��j00k�[mS�/޵^(���L���O�P ��*t�VH��QL"~/w��Ս��X���8BMα0bϹ�����ρt�($����Dm>;?��FS�]0_�ϡO��ޤ%}tf��~��4�~P�×.�D���9�ƍ���j�j.��&�P�-�Τ�e����wA7/ W�Û+!��9Ҁ�o���̐~�p��Z�^.�'<���9��I4"�d�i*3�"�ɏ�fȤ&��OȔ0<��c��Jd��������g���F�z�f���n����Li 0f^�n_�\�w�O�O�J�_�6�@6� �z��;�����9��(�8�No#X���c�p3�P,^���LO�~�F���[��ᵹ@����[8�aa8,/�!A���%V6p��T�>D��1���<�,2�)퀻����@�e�(�AqD#U˄p��L����l�l7��Q�#'�t�ֱy���4�뢅���F��E��](��X�G5���P���᫣�L��"��&y$��'o�8e��y��/XB�j31k�x�03��ǘ��B��\4���ׄ4� �q�\����v묾�M�,8!��1�
%��5u[,����R�`��5&r��a����i-<��Ѓ$���K����n@�򎫑�L��0T�A��hj��r�=�0��� ����s�3���$a�0�����c+�Dl�Qt��.�z�Q�S�22����>@mYL�4�,�`���5E��а�QĹ���8�ϸ߮.w���br6���<��'_}��v��|ܵW.�/�7�:X������<9�;�FH'0�t�۷z�,����"SԬ�$({��Ǐ�g�
i�HO�%�����4�k�O�-���aK�j�\��Ѧ���/�כ�68��~���;J�9qA��J��3�J�A�$��2"Ǫϓ�{E�zH��	�kŐ=Q)��O�j���K�(�{���9��*�Ǟ2����~��N+�q���9�e�~���i�c�M�X���2|���[{[Oa��VӬo˻^�f�,�<ו�D��>XF�l�����[�)ei�P�+ר54L���9�]�Ò�2u�����^��]�ȒK]�`g��39�#@�d��~c����kC���&����?��)�$�T�%M�5���7��y�g�A��m�3���J��2̇7�0L9yP=���6�c@��	��#��!Z�=�krc)KT��~�9G./s�A�澐���M�Cddk�W+��5i�?Z6��y�/Tj�i�e[%Yd�:Џ'�b~�Y$�c�+��E��y�A�w��T�$y
`�p?�VTڬz�1O�W�~ᦜ� ������4�Z�g��Ģ����7�P�ԯ�P ��	��&�a�Aɣ���dh��0�)IUk�3O��כ9'�=D��݇P���SK�=��L/��D#*U�!�`_�bz4���}iӳ��
�d��R���6	;�9�5u�XT$��]v�A��VާZ�2iL�$I�7{n&�Y|��qA=��W���H>�{=��a�ԣx/�D��F>,$��C���Y��������s�hl�E�2���)s�����͗��s�2�@�NG|�Н�!���a#"�G�me���JΤ��[x5Pzґ�_p,c�pt��^t��
`�B�^�^]%1�2j�������j���<���ĉGj0O��1\.E�x�M�0�ܚ��^�>��v��2|l���s�OWe�Gؖ�mX|��Y�ڭ^c1H�
ݳQ|��y�����l�ЫE��c�3s>P<��j�s�~x���0��]��t��0���D����U���J�ao� �:��~�i������#E�;VP�6��zZ˕J��!����>�J/��k �[����6�Ye"�;/�!��XVC*U颴w`����� �p(t�{_&?��?p)�)���r�ӏR3�u�Q� b�B!X�Z��M���-؀�
�c9�"�/8h���sRc뾜P��͜3lӶ����2ׄ䄗(��}��N|��7[��ŻU�Z�:��ޮ�*�V�}�<�����cF�;'�5?�� %�d�6�5���D$��o�s��2'���.5
2��']���o����u��.J�����W�������6�(��FM�i��4b�X�B�ޮZ}+#C?�|��S-�o/�9��w���Q;8jZ�=k̀��o]C�.�U�+X���>�y��6��H��m�UM��h�r�[X�J ��{h?O6�/��)߯��1���!9� *������_����|4���It&�������^��`��M�L��K���T��R[�qVY�9�;���7ad�I�LQgS-�+*����VVONFi�ʘ�!P�ξ�j�[>2�ڇ�5^D/f��� �<�PM���.�U�[\���)�lZ�%$[�2���&���vkک�Q�H}Ǎ	}�~U��7���n�J�m��n.��?���e^�6p��B�������],��b�B�Hт�M�M.� {�pYC�N���!w�P[{�n�CP��
�6�d��p��8�2�8��"-%7�q����U���t��mhȈ�zu9�a���<��p�N�@W����GK{��zS�R9��W���.��KO��S3�{��գ`^����/�PPˁ5�Y-'���u���t��n��|���A����n����N\w�y����#����n�e��	�'d�řy�>�Z��H.�D���Xn�g�����
ʕ�;`�e��}�24�7c -G�cWX�{Q��D��4�3HOw"7�}��W��^�Q��Vä���ep�+k�� �N����1����d�0�<� �Q[i��"	�fD6?;�y�<�����Y	!��L^�����ô�;�\� ǜsy��U&�������z ¾�k�A_�h��OK��on���q����Gug�P�@�ҕ{�s�7hNna��x/���BH:�02�m���xI]�GM�s�4���:��J)��G�V��E�-������`Z|�$3p�iw ������=��TI&�vӈ=���C����"L�[��>-¡����]�Cp�k�IF�d(Mʲ8��ihk���s�����?Q<����r�B��5��:?�a�U�D�O�}</ָ~��R俠�]a���v���н�L���g.J6p�(��������3R2�6N�#�pL,Q���a��ߧA2�����CE�y��FTǷ��?�KNIK�Y�9F?!��hM��G�9���:P��;��W���]O��FUG�� '&�~@��G��M:a���nE��Q�j]�gL��&�S��HTzU�}�!B�ei��P"0p����I��Ҷ�^e�b�a��@& �+�i�"���j8V�����g[[X�����4�L�nv��2�Y� h2|Y�+�1"d>-7SP�%p�������A�*yl��XH�n��F�. �g*�iH����~����� ��3��������Ny�^�ؿ��8F����7�	��(�@�!Pa�����gJ²�p���ց�1-/�~6�g˞^�	(��=h���ע�+RV���l�$��x1��m��m-�`�Ϟ����x�y��fAt���M���HX���C�����"�<N�6�Lq/�/��wd}B���F�W���u�l��,��`�`�=�����aO�C��u�b�ם�\z'�at��C���	�x��r�)��A>G����cE�����Z4��]�;��{8�l�fV�*+�	��}V+?ѕj�}��߆�Lu���}^����݃�1]^U�_RkڇP&ג	A�f�$�٭V�;�b+Bq k�v#��NH���!��U�����ASȐ!�C��،��؏�Iͨ!sܛb
�=^T�e�6�a��I��/(VĖ)��=�Z�Ȥ�e<(8h:��/MN/�����}��SE�S�B��͋�5�yx�+``GR� 	���o?�Ik����$%C���]����-�L"�����*�m'�L� +��t�1n'�|�R6�6�;�Nr�5��١�v_"��*�9�CP�3���	����71����ǽ�1��%q�["jqc��%��;
�]�e�h�`"�ë��;���m!Er<����Te���0`�<m]R(�[Z�׿�n���&�����@7�������R��=�P����i>��>�C{M��s�5H�[�¹��o*����-S�nP�č�sP�}�,�fN��Y��g�oOѐ�w� �X~<IG=C�Y��K��9����2�!I��+b���H�����;`Ֆ]C~ڌPo���f�G�ȑ�됗2+u�U��*Y1��Q��-�LC<�ބ�Ծ���oXb�R;}=Fl��3����H�ΠTE����:N �K�^C�3KB����mWm3��'M��'��.�U��Z��N�h��:73�A����G�1��q����G�K|�w����&�j����x��j���n*,2EUN�K ��Pk�$�7s��oEv�@l�}���[x=Fs��2`�c_�{�3���X6���R�hx��m�O���̤�3?��su�tm^&�$�ΰ��T�����3��(���u`lWT��1j��q�/92�F�a;��b|�s�������[NP�0����0�FV*$4\l�XH�#��/��� �q��rG<�g�Hx�phc2������x��Kz���ٹj���t�b�'*�H
�C7z�~W�F�ol0�9ܦu$�d��˞#�K)�=5����'��4�4(�f���wjj� ��k?W��)y�n��^�3t�1e2�t�H������D;���u��T��A��*�7|�+����6dZ�?����l��썦��!�*�1���cy$�tyu� �ĩ�݈�C<]�)�����毄����H2���+����g��
��X�ӵ�@7�r2��fX���XɁ��oYT�^o��;å��*��2¦4d��X�n6�l��f�\a����J�˝�`"�����ͧ�����qi�{�����pD,jtb����U^7m7X��ǅ@w&�b0����u��9	��x�����݋o����H>�Z��TM�8P1R�R{�6O��$��U�-�}���X�}s"�nc�m���X���ەzS����	ef�x8��Jן�g���zi���~�{mg]KVTx�=I ������ب���W?�����9�C��Ѿg4�AN���=�"y����8�q�]N�nV����F%�.�0 ��]���1�2���V(��P|g��Q���u�-��'f}�_"XTҍ�H?�m��3�!I����ٵ%�c�P���k���J��J��M�"�R6"}t[��[�Si�c���/�V>�%n4�����/��u�[d6�s�A{�*a��%h�r��X�����e_��39����uE�t���	��΁�Ws[;�i�M�	�����d���C��+S�e!�����3��f>��+���W���U������:�],I��g������e0�d��/���V�-2���j���Ȯ�?!3�ޯ�m?�0�Dή��"K�?�̥$M���,���'I��-�(f�ˆB�����d���˸�0�
�H�������iQ�����W4
L�#�&͒�l�&T���N�>S���9t��L<]��'�]�@��8H���C����Ɨ��弡 �dB[Y#!qU�>M����e&��N�,�u���%�l�4��~�`&z�[�}�ϫ�f�W'oy���1#=�Dدk�.q�(��3Z�3�_~x�?����RsǆD�	��Bp��EpO��F���3-�,컂��G�4�B�nG'��+���xV�����}�&?+�,%2:r��|�s�j��=Z1��3�2I�_�{d��4N��h%h%(G����׋�Dߪ�w��~<�B�૿K'@���M$���~~=,V�X�Z$#�����(��Ά�í�w�Ǿ�#��ѩ:N�-M�L\�Nf|����J�W���P��jpe����CZmI>��֢1�G�9���y�9��#I����O(ތ���I�ٰ��Ǿ~��.~�]�5���9Pkl50P�w�|Ud5Rq�jP��:���8#�/��5�����$�"^��	�>:��X�4`��<���X����)&vS
�x0��@aM��:U���F�=U�^?{��lk���^b��Y�Z�G�h@�)Oo�>e�Q{�#%Ȓ���1��b<���\�̮��0����d�$�(�$�ԕ�������A�����"3������k��R1ҵ&��:�; ��l9C�O�kʵ/�K_�45Qc����x ������7�RISI�~�U�=���t�!���۳N]�F��vǌ	�0�Dfթ4a�u �n��{t�t���O<�����,z�'�<hS �]�7yg8uPi�o�v~��N2��l˽��e8,���#f�Q*�iv^�Rљ߯�H°&���KDSċ'�iG�|���P�"����;){����dfn?�n���s��n�u�SA�U��kV�=1x����љ7e���S6�׾�Kk��^������䶬pꏦ)��2#j[��H�j��#bxD�;�84�6�f�h���6���$p��t
��p���;��}ih��Y�1;Ѕ�آ���a�|KU2�T�qzt�.pY�(��,�"U�"OHp2�~<S��X*K��0�H�ȿ�U�5z��L���(-�긠��;�m⌚t��X�95�Lw]O�j8���̂�>���ϣ�8Q@�a�:�l�t�j���]���g˞�f�$�2|��տR�sL�N@ȟ���Pju�M����T��H�I�������Y��4�'v?b� fQȚ9u�eD�0i��!�~L����z�
ˈı�/�t`����p�E����J���yN`���.���5�����}�Z�p�Ro-���>!�^ܜ_N��g�G�	�1s	ܗ8a��n�J��hHq&\_Uyo���l����9�����Ռ�K�|�w����vjǁ$\�Ioj�|�y~	�Q{x<-��Ev�$g �P ��̄�$a-�Sl���q�S6H0�Iw9MB���L�sv"��6Y?�4��]R�m!l�Tm�Q����n�d��i�ל�G$+�@�|�^R0�p�)���i���Jr-`;�ţ��r�ȫ��2'gs�E^Ѕ�� �2�R��m6��r�"�w�sS�����%�<_G��y1�Y(o�UO){�����ڼ3����`�^�|��/��2ݽ�α�^�w�:�r���p�>\hI�,��睊1�L�{Vk�7G���N4�N:с�z�<Ʒa�� �5~����r5�.���j�"�i``��^Cv�FkK����яu% WG����y����_�a�����"��d���l*�@N�FVdT?��W�0W��`<UIы/u�ᓥ�'�Nq[��V�dK�G�O}�`I����6����az��\����Q�ʕ���j��g7�B��{��+�8"(Y1=�$o^,���l������`��u|��U��I�[�R���`��a^��	k����=A/��a-<������������@��9�LT��e1�U4�d��ȟ�IK&6���֕)6*�#��߃��M��u-e��_3f��o��qʐL�|'�r���M���ǫh���e�O��o}�����J��+���L�v��&<Ĝ�.i4~^D�ԅ��cf�#a2���x(eO�oM�A~��>��̜?�@� ۻ�-�v���E��7�;3�N�a�,�3�?�-�7YV��Q��+H�yŋ��T���-�e�1����,=4Smgn;������
6����z�Ůf�c/��J� Hc+�ӑJ��F�] �����EЀ�9�����I���&�~+�w������Q��
b��Y�8 -T�����;ڸ�~ ��N�T����.x�}U��Q1,���4)|�$�����\w2K���X
�/��}�L ��&���E�+Q��/T�<�_MdD�WB3�q �52��/���$��d�U:��>�*n�`=�֥�(+�a[77g�m���]��_k�*�E�Yƣ�ied�Igx���`����vj𭙎����*�se�<��4+
�|�ߙ��8�.�B��sAu�ɤZ�r,�����?�
S�"�_�:�z� ���Z�8y�H�������"qi���u18P)c})�c�A~��q�sa�	5�"��c�#˹��B|���D �4��;Y8����o]3�N�i"�5-R�F�a�<��U9u������t�B"$�����tuh�';���H,�UqE���6�%�������%sh]"���a���(��@ޤ��%�mG��5�T#0�tS��|��xD=�]ޞr6�7_Kgh�[�6�]�l�q�؇�{��_n#��!�M߬�323+C�����y${	\}J����d���9տ��Xg�'��<H-T���ʠ�5�^�:�{�k`<]�~\��"�L6��PRA���t��!�wU����t�+3bX���:f���`	�~�A]��1q���������.���?w�Y�<�����g��]�#�S�G�G�cy�t�Hܳk�t@7�tVI[����� tG t��l�v��`"@(�L�$�4��\��7ϔ>�\e���Η�LA��:���͸��)�h��j���~Qص�.��y�v�o�fp�u���>���1:�	||�5e �ݳ�2L)R�RŒw��c�2�T��-K$g[z\%��׭�s�0>��"o��|h:��~d|:u��`��o�o+\�o�r�}o�9�Ox6��Mi`�|P�8��0".��H¯g�%���^����ڧ�+��r��,��������o��n����ֆ��h�D���;h/��,pwkB^+��&�|I��([��nz"�il��&ᇾ�!ȫ�=ΡR؞���gO9̎�$����ƭo�=�f�_�*t���{R$�)þ�.9D�`�s��ȋ���p" [���(%k���y;+���}_�Tm���w`U}E�,VK�� �'w6	;�q���_~F� Ĳ?���|������ě�\�Ձ5�r,���j���φL�Ԁ91^m�ôub���z�Z�ܥEʃ�ʁŀ[��E�r���kO@��&	���G-��	з���k�Q��PZ�f�l 3�M�A
�LIT��%�~��Y[�oS��t�^(-K��g}��j�1)@���Y�B�	�Fµ6j�� ��Dn����ުV�o	���݂��yL��wQ�q�H�ZT=��������	{����:�L��:�?��>믕;�TT�B�amW�X���/�a%y��+�OA���h��!,����v���-�ѡ��T��7j��n
?��y��$O#51�x��u�Hc4�-�����R�Y�����Ķ�7��h���\ѡp>@�#?R}�~�.k�!��k� ��P��Z����N�/�� �H'�Զ%h�`���a9O�er2���VV������L�~B�|-�z��Rɸ��了�F�!aY*�
��ӣ�&�}��=�vjz�(o��� 9?z��7���O�4{���C F����NaP�O��kM�RY�1��Z�\Ѡ�y\�;�W��٥jYm[ݢ�CI��iM�r�q�R�<+VEX�M��]{�e���.r�ϝ�/��w���q��ŋ�4�M+ōP�Э�7w�
R������B��>��i��p�g���o�(�D�t��Tl%'{��8}���"�S 
��hDuT�L�PT��,�+��j��(ϰ�g��9��%�2�E���
|�JNn���%�����kŮ�ؾ�é��)\0�ʦ�Ì��[^����R�GXg7C����Rf��^�c����P����z�03���I�ig6�!+�-g����'�����В.s�dM����8>}f�\��j٢Y:}�U��v���!�{H��n,aڈH�fk��$��9�}= tNa���͆U���ٔp��8�6?���\�����������WI��{�ö��R	��62��n�#���$�����2���ߑD�����5zO��MGC'���-|abHTݐ!g\��Ɖ��7��r'*�ŗ�,�@�HЗIX�_$��[�ޖW �HJ@z�#���n�-
��c�'(>���51G�W��~��ﬨ�oy�J]l��=�@o��UCP$�:�4M~j\�����j�o 5���4[%
"�h�R�Wf/2��:�����k���xBJ�ˑ9�Y��I}9���ߵk�Nݿ!{��d��;���0$�j���3jnty�X��0�ZIȭ�b52K�>��p��}M�P-�pei�;0�x�z��ƫ��U~�j�Hr8ի8J#r�t�Y�##�T���м�B��y��������<՝4�
��_Ԓd>��̆�_7�XJ�߸�HR�\���\"�/,��;0�j�?�|@Up������A���b3e7ǁ����9�l�;�� !3�̷*��)��x�_���l;6�or�L$�Ag8��K@���
T�O$:8���E�H�yB�	��iu���,�#�i��G�B~9)��?��҂��07��ٺ�f���Ob~0x�%�&�w�X���Xd˧�����8>NqQHP��&�����q�Q\����xs�)�I���� Q��r�m\@踬r��ƣ�t̋�����a�n�O0�3�)�r�h�'zIq|џ��|���ˣ���K������z�����4��}?f�r��X�OH)��q��̓8g�	�g!���m�'j2#�x�MG�=׷�ۅ�n�Ѽx���'ES:a��u?�k��F�h�v7}B�X�������S��$��6�ۑ�ܴN��}��K�p	�|���p$+�̣!����Wt|�zm�j@���`3�<�}�pN�Z�MY��I)d)u�\d4)("���ӈ͒���?���Q/"[��g�y��R�yS�S:.���
�E���Z<^x]�g�>�,�m ��(4[����Ŗ	o��S�z��z�<���ޜT]�=��/�'|�ӧ�ǳ���������orS�'f���Z\��D����
QZ{ll84hS��	l~ƀ�S
����R��+���mq�%ݨ�����AhZl��}0a�lM���-o`�P�n!��z9?�fd~�b���݀6];�J0E �����WH�|�|�U?��F���3y�}7H�27���̗3qr�P�������%�{f��I���z������R*��j��e�!���D��\���+Z�#�	�?�
�������҂3���Y2���5B�Rf}k��¬[�T�96�����.�&g��Җ��L����7A��3NyI_�=� �ȮmD\}B�l�dq[��2l��A &q��#6ϕѳ���þT�{�a�2�/��s���,���q��Q��]�tU�$̠f�O88�0�m���RP��W`�Mh8)��}|��Oq���Z,�=Y���G�Y�$A��>^�9�TH���� n��ƛ����M|̓ 	,w��}�߭Gn@D"� .�Z	NY�^Ǫ�ֹ�<�Hi��/� i��G͢%���,CG�Uy�:�]"\�)H)��Dr���4u��?�%�(�Ā����afĴX��ӵ1y���wM&L���/#L����J}"��ړ�Z)Ҧ}�~pe�{���eTTwI����0I��� ��#ypF!�k`4���i��Ny�e4�*�6�eG:�ʌ�t����|����Xm�E��pICu�[���F��B��<�)�NMk�E����'�ۛ�G�U ���]6�W���\O�`-$op�BQ�u���Y3	�8!>��h<<���]�회8P}W�4#	i���`T%�<�)^�G� �O"?��;(�{�H>��N]+��:>�ys��1�Țه�._j:�CK�,5���>��H�k%�L���E�G��~���S(�_d�N�"(b&Q� Y����3�B�X��W�d�і�U�����m���u���ٞ�����(�X��W-6���6��ծ���a3������	vv�
�T�vP�����$z��3��ƹ�c/u�\K+a_��M��ω��b!�g4|q"j1��Ƹ�+�hQ��5�͐����A�a��}���I��R	��*��՚@Q�
�-Nm�x}��=�$5�F�Gj�KV{�`�����@�g?���T�N�c���;���	�&���$����Ȏ��< ���B�Y����_�k�nBWA#�7W·��Ǆ�C*SDޕ�	��,8P��#�?�C���a֗m>OC��M�DRC��!X�/�]�a�C���'�Zk�\��X���O�,�+֗�\�D�ԁ�I (*P�ִ��g!�f+�}���	��Df��Ý~�`�E��'[zaP�A�EV��v2�hh�NX ۞�/�זN< '0��փ
J?/�������&�=���gԈg�8�Yfޣ?�t�T�2$��ʈ�f���1�i���@��?�'���H���j�ԯ�0��L�E�by�(�L n��ZN�?�Xs+��Υ8�\��-�6��j�O񡾳a$��F�]�=�w튻νO<�x����ͻ�����w�;�jR��OL���X�!M�*�5F�Ty"��<%�n>����ء�׏���f�R�.�E�z�t��c�j[�z<��m'�:�h4/F�y!t#��&��]	O,�XlJM+���NVak�-;��s�#��ř�{�,w�"�Hl��^oɜ�%F�pC���J[p��'��~P�	f�S�*�[��h� ���K���q�����s�_�ei;^{�x�������f���2���%��b��A�L���4qt�]o�c�}��4��0�s����_H���,8F���,v�΅��N���-���T�����.�6��7_aR�Z�]���:��/Kg3��S:�6��t���A-���n��:�N�k��ɒ
�����D����T&�8����0��]9�m��{t�rq�������4��3�B+�!�$�NQB��-��p7�� �^��sC�e�n�j������+Kd���fVUSLe�&x.�l����Ho�e²�'�|�51g;���^n�y����!��9'�0�S��ٟ($��tЃ},/�|%�1GD}�g��B���ےhE�(%z��:�[���ɽ4��%�g/�b�2A���~�~B�KT���'���{�U��Q0{�j{'�7m��
���0Y��֚&�����m;SxX-ߦ��͂9b����u^TQ�Y}�f!\-�q���%/tw!4�����:#&,�|�[��?��S�xt��#f�DN2�)@�!To�fD%��G�`i�k�[�{�d ?K������m��v{QWCI��Lh�N@��\ҏ��?%`n]N��2T��ji'#(Gto���*��?u7���aU]�oi%�/�ā��i�S�2�g�'N����aPx�"�8���/"M@��x~OQ�'���O|��l�#�_c�^h��={�ֲ���Ʈ��3����팘��s�?1����9uV�u�-[��x"W!��6�I[�:�z�Wb�����K�ݰ2+��V`���1d����E
}YPUo�WoK���ϱ�.j Fh6##�f�f:� �W�:�_��nw�kP����Uc�/�Y�\���ĪZ�ǉ���N�����t;�0jD|F ���A��9Y�X�{k�Y��ﵰȶ7�F�?6����dR�K����R2�6�Sϊ�gͷ'�4B�U�<�B�	(���Y�� �{_��w�d$|/�W�]�̥�iid��pl .hvfN�ń�}�bZ}���o%�����-���7��Q��`�f�b5���.����M4u�1�kgZ����WB�9�Δ6L~��ڔA���Bv"X���؅"ߴp��W4�N�|܎��5` ?�������tgw���a7��Z�8T�A��;�����������ӒG�(\��V�*�������d�>�]��� ϫ�I���c�?���t����0�W��|F�9RU��
u٭,�;���J����t����ΘV��c+��ғ�:&pX%��7����P�%_zc,&�{O��ؼ�O8�m�~��A����o8&�h��.��c.vp�Fڽ��_,���E$���*� ���/��>j5y�VoN�l ��n��j�y������hl�b/*���H��(����Sa���m�-Ww#������V��^���!�VE19�����L�?�Y�x#�����d.MW]�v�v��킳Q~{&���\A��oݸe0�"ܭ�;K��%�}BF�wꉏ%��:�S&��N._�N��b��'��K#Iw�c�=���24ಷT�9���#�+d]�8\_�FU���y�:$W��p��n7�ȭ:����Ә�z��yXҸ��K�W̖�%k�0�,`�{8��A}N��)�{�ơ��/�nhX{B��}� �-w��2�^��bv�����r�ShXFy~tE����Z��bw\i�H�0L��ox.�3�qҋW(\�GfI=2�	�4%��Ny�Ae�\���I:�|Wd�p%`{*��D~�=�T�c@	�II�ji���H�a��T�L�u�8�{�5j�u��y����H(5���Q�	y�	}�+�?�U�i����� ^��S���w?��w��	�#�}��B�5��IUwΒ�1|@
�3�zRG?�P�s2����-�$�.��^��:�~����F�(���Ѧ���zس;�	����5ў-*E&�ꓭ���ʏ���4P�O�?�y�^k�Z��ҥ5m�W�?�Ã�T��\vN�J�-����_�}C��][����C�w��o!K�8�{�3;��z�J��mj�]<cS�0n� ���h�.r R"W�.Ej�m�ѕ�O"������]���Ewن��*���M>��Kj���li���(x��ͬ�]`�(R�h�Ak5L�l'����I�p:�@��!񨹨֤)d��t(�JIܟ�(;sJg� ���B��n�oe�SؾG�*x�i�潉�����ʖ��%ɟ4/C×obe���Āk>�Z���` �l(�<uzȲ����m�c�_O��6��ę=n�<W<�2on$���I��It���K���v_��d'|&��p"Rn��"ԹC���Q��-�����Dr󰵝�����,�?��-:��,���g�/��ՊR>������7�x��l�ľ�T�fҏ��~��d�|�;�a�	�S u���WN�g?p�a	���}>!�5]~�7[�g�2}�a��J�n
z�઻`U��b�p��EŃ+G�������߈Ī��!�+H�2�1k����N\�����3mki؛�IE{��R�
?���:�!pg�IXdK�{֫^�Ͷ���G�:A�M�L$W ���)�M�{��W�=�.�;IqPB��Q&��|�d����C	�����Z:Ię�C������<�7��:v��^[	$��Ȗ�M����1�bR��Z;�>]�EDk�Z�'���zVbH(�
f�U0�M\��)�S��6'�ײ��l�}���O��E��.� )5Ϣ�r��Y�Ld$��S�&f�xs;�"]�K)w�S��4�c*���(|gT�z+a��s��a�Х�A�Z���VC~I�#Fs,������o��1�z��n;Y�K�/h�y^I����_6�Ȫt����}��Q��4��|��ŬT��tiUT5�^�ohUī:ر/�`r�Ka�D��s�l�a9�~���	0/�������5v|M�"Ԫ����5+m6{����~��Ψ��HQ�h��Q�|�v	G��a����[��="��}�l�1��m��P@��:�Z�ʠ�;H�z�ֹ�P�w��"���/��ۉ	�{:vX?&~��{��?[񖔅����E��+ /����a C��"����?�H�}`����>�Z��/V��2v��+K�ԙ���_���2����x:"��J���`"|��s@��Hw�ٙ�is 폞�[�N���`�_�/��TOM0_{�l�(��r *fܷ�~� ;&e��f!`���^Q3��Ux|����0Ѐ{�i1t%%�Iwo����7��� �����PΚ}�B��&����j�X!��XN��=_d�v�>Іn,uR2���v�.��+B���%���霘�8p���n�E�]�����
n9�51F��p���H�dM�����*���[��f _(��������둏�cJ�������TR9"�pu��Ehv�q�P�tz��$oΜ�eG_�s�g8��'���nlv�]�m�2
�|��� ��&MV٢�6�o�`��0D=�c�K��k?k�Y	;1��]k��PL��"����ӷ���@�q�0Ѡ� �:���1�����"x�0;^�+�RX-"�#�T��\L<+�MoL�Q7\<ڭ���))���mҥC���
;Hx L���{q���<�H�d�w����j�6�t��u��t��3[�W2G��Pk�5�Y�`��_��,��+5.�h�"�Y������9F!U��&�=�Z;�K9`�ҍ�CЋ2��t��:�v�N�9��r�~m��}s�1 8�T�eU�I3��tv-�*���e���Q!J���ל�b�v���A�ְ�!$!�˩W���_:��Ts����N�Ǟ�x�\͔�j��.�"�h5@�BI���E5"LHl��9���~LQ���t"�E7U.$�MԟeNK�[6��=�A�,u�BH�y�X�r�>�6�#�iDϯ�\Lf3��"_�z�p0R�:�m����8^�gR���8W���?6 �!̙=�D�!~�b�	�W�X�t�#"s�x���:MDsi�'��5��QtV�$z��jk���}���q��d�iƸ<�E9�و)(��Fo(e�}SJ���r�8A��i������^���Ԕ΀�_��, ���'r�Q�=�!�����ޅ� *{��XNZS�?SC�mԧR�+T��	 }�t��6����'5р�G?\}����@�?������k��@F�x�@L5?&5��$3;v������n��4�6�Ǥ�]��Jx�i�3D��	�M#�kY:�YDE���&9~�cέM0T���l	1�O�v ��f,�ٚ5�0�r)N���֥=�B~C E�|��C�hw�����|+P��ᆺ���}��b�>�5�7âR2�}�U!
��V1/��L���ה��
ԃ�t~�}�'����D����Y0�&�"Po3��U^���CG� �q�?�m��M��!��H�-)5:�wEIT���e������Gv&��33�C!��:J��6覾�>d�1���U����"��h�s�4������� �>��4~K��&�Ŋ���8A)]�WN��lî#C1UP~p�z�.Pz: 9t�� ;��@XM^�!�1,�8���x��i�?- s>��7�4qq�RǭT�P;e����W�"KU���������b������~�_ ^X�r��k�1����2)�����o�m�H��v�S�^��9��s�8��&��ttj|��_���ך��[������xN��[��X�v�v������S��)4����0�8t���h��#�@'��]dˬh��9���}�@�
�� �Xd^"�<C��{��v�Q��TG}�ɼ��ǁZo���΀����t�&�7o�<���|]�m�m��ǶVp5x��#�d8a{�8dGOȢn�_��<l�e��1
�L�&2��\��Wj2ɚ�ƽ�J4����$><-$s�gl�@�驒�4[�]��uh�D���71u"N7�wx&�cbTG�,F���6�]C����go^zh��Nvi��av�ﴣ�/�[�Ɩ�K������w���Tq!]�-�*N=�c]�gE�Z�����!�Kq��[ٵ���ր�yS���@�J\��n�)��zz���֯�4eщ��rT��7�L�)M�TT���@�J�Bi�����կ�t'6����MJT�=���lơ$�ckRjyd��j;��0��!�4LF�),(�f���*�G����&�����%U:QWkȽF���~'�a�
S���u��5j\,+��uh˖�sB�Uc�@�G?�3*��~,lm\<���=M���`��.6i��!�@��ŗbhuçf���_�̽��d Nۻ�9�c=�x�����r���r�"�Kpk�;��K��Ѥ֌0F��x�s-��?��� �t/bH����(�fϋ�**�ھBri ��;N�;bY��Vƌ��4��@�S�}�s�μ�h!t��Fi���
���-~�j3}$G\��W�_
�@�q,}�Д��e�h,�:h�=�°��v!�*f0��Q+G�uS�ԝ����"`a�k���2�����ң�nC��]Lt��2�vs-�
aܱ� IXT�-w���Ζ{\w�Y�p	��c��*����\!��E�'C��&"|��x����1�� ��E=�z��)<=�lø��� ?)���S�i}N����w�
]�����*��kt��h����RL��8t-��v��@�o1���Q�|���Wo�9�D&�F<uI���h�-3}JN�^T�Ue&{`&�j��$Pa�F��Q�Qu��M*m��l�9�~R-�E��D:/}��
'd;s��\��0�<���8�:{�б���*"I�qJ�q��p�����H��E.�ń�M���MТ7�ު���u��v@�H(I�6�Y��.0�0*VD�t�\���CF�L�J��/�7�E%�b��P��ƃo��~�2������l4��4�~� �]�C��;O���݈ԺF?<�En1ȎHAA:����J$w̠��s��[r��Y�1���(%���o�#�u��E'�X�����x<�#g$�P����M�w�]P�wDY�^�B����3#xQ��^��k��t�����0![�)�"ITK���,������ѝ��#��.�E����t��-�Z��_o=�����+�"?m��V��4Z''��E5>	�#�J`�	��a��:���0����|�����{4�T=�E��3*�?����cܦ��@�KQ�g�V`��ǿ&g9=�Ic��c��w�gwbʃ$=�\���K޲�8����ɴ"�r:b_Br!�D����ً���GيX���%&�0�^JȷW��$��F���� \�|�/pS��Qw}>_#��W��ɿh!zmK����/u�`K��
��!��VS��=
3�%#�1=3D�f�op-N�|0{�Ng�f��t�=�����*B*OH�C�AQnM8��=��힥'�[ ��㓋4(�8�!	����-#��|��d|:�&^�x���?�Eb�� �|z&�7u����4�PH`�mȠh(%�L�U)�l�m�������	Y�DǴd��3Dx�!y�Ҋ�2y���v�\C��̓�,�6Ta����s��|1 l��gK��|�kE.��e'��tm��c�Xr�_���Z�ӽ��r��·׊�Z!��ʓ���8�� M�.5wW�;eN�M�����U��0��P�#�-)dT���'?��N���R��T	Ui�0YKǙ_����� ����O����g�ǯ�a7�/�����&ۉ4W��՜V�2�*��d���ƈ�ax���E�Q��⺄����W�&�?4����B�)���F����ɺ����M�Pk\N�"���,�'�R�g�5D*26�-��8��h�1��UY��%�%5~�m5�l�Bϸ���tt�bՅ�C�d��+*�l�ת��b�4 =:�vos����@�.�%.��P��䮳�a����r���o����a�y.�	��5�ߋ1�	i.v��>t���8���!�uA����d�%�bx�Ug�N R��6m��q��O�<���M�־��I�J�\X�c㇡�?ې�
6���� M����VgI�l�,I�L���.�9j��"���ͺ���4���II#@|�y#n�-f�����`G]r"���^�/�mڽݹZ��Ͷxd�P�����U��ulj����o(�����(����(��c�Nwq���r3����UT��.���6��qĎ��u)�������G��!1;�6j��F\/):�ǕC�7�� Q\�*��F�G��V��Ȱg�ef�fzX�Oyj��\�I�:�w�1�m�_]���۫�B�8G��Mhҡ�T�8�(��e|���s��������d�+�U�u#i0����q��^3l� �s��-q������J�����N��:f���t6�����M������)�\����\�QI�x��E��_�y��v�Q��X�J@�S�!�}/�+�q:UNj��������{�q��BM'�����ôEI����N�N��׫J���~�[ B�6�R�n�&���G�w�[X~y��b��
��Vd��Z�_�G�}1�$�-(ф���umh�b�(��EqPS!�FI�%��{���Ȟ�׸5�l#����%}X�e߯�&G��W���
W: �[��Ӿ�䥴��#���:d?�П)po�iI�?��W�*��s��TF4掵��O���_֦r	,����\�	r�ʸTeAmyUi[�u�����q��h�M��Q����-�	&H�¨��O�szdmU�"+��L�4?E-��m[&�YtHT�>*��6�8�s
���ˆ��HߜL�$�Y�Tܚ�y�b Jbu����i���r4�9(Dw4��aO����ހu۩�qǋ9H�ⷶ<K��1*%wh`)(�گ%ۇQ꽖��,�ۭ���V)������|���y>�A�f��H
 gB���0ܙ�=��c� o�uOv/u����p��q�U�,��$��)5�V��2�A��r��헸Shh$���F������|�/[�p~����T����ug��<F�>�����b�oR��==u�O�F�U��f���y,�w��1a�񲯕��i�J�kC!�PzWee���'m�#�K���+ �Z�,���N9��X��"�S��������GF�s�=���%���'r"ڦ'^T�(�[E5=K=ْ�d{Z��C�1����gP�#�m&���ҰWl������N�J�֚�<�����%䥮�9�wy7� �*Tׁ43hڭ;���K�vI�M+�A䊕?���?l����}�$׍��V:�����W(LYj��)�x����Ju�;4ɱ�����@���6	�j�%��0�i�	��z�O3��zv�h��8������`�I[�D�PS)�X�GF,$|A{<6�vЙn��jq��q��T#�v�z��L��F���sJާ's4ˢ��\������ �� ����~[��z���O�����\���ѳ�pq������+���8�}ǋ��Ae+8/0Q-��I#9��S&GWx��!4�ֲ�)���6
a�AO6mA|֔���������)"�#	Ͽ��\������V����D.����6����:�(��݅k�68�9m+�i�Z3d�񭵏�(+<����A�8���D��,HK�/§�+]He���Q�={�&�k�a��C�U��QB�b���B���T:��ʑ�%�"�{��6����,�|a�د���P�X�籁.?��ZQK���gRܰ�j������r@��lAړ�<��kᜪ�������,N�P|�d"+��zd���꾬\�-���5AUq���B-�1D8$�4��dBC��5g��"g���r��i�������3�QQvY�ʠS��g����@Dk^ ־C#���Gd����Ԏ���,'u��-r���0��P�^��d`YQ<�M~�2����r��8@��žBI�ѷ:�	ٖ����'ů����U�7���Rr��g���YV7IU~��g�9�+V��6G��>Z�=�y7���[�B 7V�'��4�3�n-Qϔ8�kli�͸�����{L ��MN�KV��/{Xɩ4��X(�םnP�s�'�Wԅq7�}�>O�^�t�;�c :��$�%�Wì�,��Z+����bJ�˩�R��|���h>Z�tl�
�rTC��3���pW5(�G�2HL���x:���<2'�y��1�}�y�7ɜ�|�K�~t���&R��}%3x�Л�W�0Vb�X@��%n����)��:e��~74s�B�������y@�׻�RcK�>�p�Z��7�`]�x�;ukĽ����� r���켴�^�}O�Z��j�3ż`P����X`��ѓzSb�?V�n8>pn�
�#�.a��s��������떢Ia�j�Iu9��W?��-񒘭��?�fyd�]g-w��������S[F����D��4D�����.&E��u�8����Ai��~P���L2ȣ@�[K)�â�Y��<W~m|6	M���W�����_c���РW���
�Y
�0s��ƯX��-��y{lpa!A�i���p�+,����J��Qd�6�n���,6������Hpa�ٹ�},�'�؝�%�b���(�d׻������h蒆n`�ÞV�]�3��c�=��:rs���t�} �Yҗ<�צ��zИ| �'�N���nޯ���F�zёa��9�x$�g���P!ql�9VxK��6����iu��v7�*��~G�|a�-���\���4��E"��xN�d�˟�
���{W�>�H. a9��Ͻ����n0�}-̈́yq���M�����i���frlx4�U�.�[�B%pIe����Q���T����(�6���Rg�ۋ�'Bg��R��h{+��+ŏC"�X�F����v�ATM?|��%e�MAr~N� 	zUI���k�]�UCS^��Uɕs8T���G�u\���WѪ�EJ�W���k�Z"�=���o_* �/p��4�R�`�6�a$�f�.J��|�M�arI,O�O�B�\1zx���f��ʫI�OO��d�'�U�u��;+�<�-?g��9�H�zX��Tډ�F�iO��C7s8�{RKe;�®a�ܲђ�#�y��ce��>YO�A����1ϔk\��U������ř��ߎ��v����ڄj�M��D����w�f߂j�S�9���v3�t+eZ~P�8���<;�L6�>�5~�>s��;��SC��č��9��Y0=��m�fW��2���Ɖ^ r��t,�j�Fzy+#�;-����u��C(J
�ë�1�9�>���'���
fpb �l1��c�	�@T&��J�]�#j�Fpߔ?+Ξ�<�a�'��U�*+�A�3G�9@g��3�"=E9V�q�ePT>ٲ���(�u��'B��w���P@����"/$`���F�*�� y��TI=i�@��YS±v)��*�+C����J����f}����K�!l �_����w9K��-�j�ʵ u7.��XGS���Ț����P�3��F�����X������猡b�j5̷��ܦ��~x����XQW���V�F�#>�n؂���~����X�sL�`VG�O=)��b_��l�Tvr���aZ�!�OI�ƋF��5��d4͚����ᨿ�T_
E��-n�Qa��,9���]�%��;/Y�0��h.C��&���)^j� �f�\�7=�(Q����Ҙ$z�ʋM>�`Õ�;t>#�[�8���j��I�S����{�B�qj�a}�e���]9�d$��I��sfY����w�7\�*Cpn�h��5-V��('�g2���:�/�Ej��f휿XHZW0�~(a�Ӻ��ix(��S��:�;`����曩���V��<����˛��|����ӫ�<㍾���6�.3�K�ơ���/�UqE>ŵ��ֳP�j����B,��p ��m�����Pwm�B�|���2k ���񛿲���Yڞ���Ѫ�*��Ѝ�Wf O	I�"=��5�i??��~�o$��%;v�ޏ�j��R�� ��7N㹉"}��-$V�o؞��۵��I��#6�;��+U6ϟvI�?vo1I���ϋ <�%�k��Xjc��q�e@�h�z"88�����d�E7)����P��<^Ѷ�B�Y���F�S���O�7�G]��|ၸ���`��v�J�6�[��
w�Y�ZX���xtzt���Y}TBQ�8bk�P�����
�Y�5%�QO��n$��������5�`�x1BI��ߒ���vG���\����L�?�QG���u�8Qq	��#�.ew�:d9����3�g�ߘ�	�J��ja�vҕy����I=A��P♢m�t�4�+w�Tq��ά�2�SD4sL͗��D�բ:���2!)�+�:���Ҵ�N����<��VA�oJiɲ�����GG:\��]�8��B^�W�(1��̔�\[�n�[� �d]��D|��E�4==�~�O&�Qa֚��V���$���d!Y�d:S5��=��/��{�����D�Èy���Uc��?�N~ؒ
����O�
�U�V��O�"�C]߫s���n���k��e��?�g����eԪ���'$��b�5���:�7K�gF���Ѯac[�qE��뽚x�����$�B�S)��3ɇ�(	���.���x�t���q~.ABh����Y����B�\"R�lb�c�Ŗ��z���)6RT��N����o�6J'M��#�7<���Z��b��\���S���dZ4L6 ������!��#��|َ[�}^�\8��N|=�.|��
ʚ鬽��ub
e]bB�N^/���-����8j�l�Y6�{�z�� �����d>0�u|Pc�@9�t�`F�p"*�lm-���^�ƿ�?oA��T
���B	��v)\hdWf ��	](�	�x���wn�W��o�_D�F�fcڢ�@���߾�F�?�`�w#��x޹�(�@�����`�hI*���m���K�n�bR�Q�a{�� �ݧe�������d�C(��He���Yn���%��>�!�W�^��GEc�!+O�I��6�7�R��4Y+ttQEvP5��0*@|�<��֕���iXrS���"�e��/�Y�D
�O$b2�2�K�}�W����V�&!�(2S a%/-��u�M��O� O��5A��N���4��F�����q�d��^E�aF�ݰؠ�����-�N��vE��¸I' #�p�F�z��y�w�o˭�x� T:/�.	�-V�a1���j�����p��&Hټf�+xHN]{]Ґ�Ϧ����6�6{������jw%	��Fn4�k����3��x��Z��+�
UA�ha��1��R�P�Pt�/��X���<؍N�e����Έ��]�n����'E/Pl��k��K:B�m��=zsE��1�7(�"1�aK.��ݾ�.P��\���CS�+hU+���밠0#W��׶��9�x ¥ֆ�rZ(D������qa�lܻ�0A`�Zmk'�j�7�n�S���y��D��qS&���AycB C�$��:];���M��"�r5ai.���D0{*�6��r��!20ОKk-3�㮨/�DiFrQ��g�N�g�BN��J��̀�2'�)�A{(b=J��
M��ȭW��PL�2�;�����KT���gc���@Zh���L�)��%�;��nӇ�߶0���DQ7�H�Nj;�mߴ�����U��4G>{��jS��M����ҳ��bf��Y��X�u����2N��g��)3R����w�ң�-%d	������n�袑�!q�i���s�+�����F�#�l�^��y��B���`H�1��h��=�6��r�ɔ�ym�
�Bu��u�F����� ��w��#[�2f\p����?�A5����8��8��"�����6�=N��ϴܶ������C�np\�WDИ���k'�#�uYSOZ2�"��i�
)Ftfi�n�řj��2����V�E(f�49H�O���Ƒ :��Q����f��5.׳�a_�������-�ߔ{6=�\��%�ܤ�>�����b���I� ���h�{MZԐj#�Y���le��?��,z1�~�b��ɫ�qN����@�"8k��1��F ������f�C�%�R1�p�MZ��p1^���e��Ż�S�{{�=�?���{($���.J}<��=~·�D�F� �[����z|�j�%P�<G�� �y��Wvz)9ak�����I�L��s�Ent��\�#J��>@�7�C:��������Cl�v1El���b�V�7@u?����
����pb�r�@""���I�#F�nݶ�#/{ȍ*��'[�B^),��B	�� A҉��eQ��z���r�;x��{��_�ؚtc؈�c�0~_�%�y�m8b:G�B�Y�{�^P���cUAߞ��0Q��&�J��7<�ޒ縙�l�;aU�R��YG?n[8��1��Ý�UJK��y�r�f��m��TʺuI�+ߧ���'NJ�d��K9nͤi��������rvN���1	�M!H��QUk>�ܗ[�a���P������;��ȹ�-����\�W{'K�۪��G��A8K�Ŀ�1p"z�{^�y�W��<�7~�����uP���]`S~�F	��ct��qg$�F Z�T���$^ZY敵Q��r����� �#
<Kڃ�A0����~7oq�I?b��_J�+:�R\v��#=v���.��.[�a�5�`��v�	�q��)�1ohdeq�Im�x��c@y⩗� �y�Ч=;��<��A����]�/��ƿ=��_�	R����� �6�*����s������@ǫ��������̏$����.��.>M����h�tFQ5MO��s�фr��1\"�^��E��Q̹<��{���*;��ś�������S�@��dTT����B�έ����aHX����H"���̖�	|��bY�+��T���&�S�s�U|�6�6"?-�t�O#�D�V����J�㽊�l�<@h�'���&��q�(���)�ш�4v���Ւ7�,�2�%�1�57�,Z\�#����fr$�F�*���לJ*˶�=���������i����Z����{y��۴W��gQ7Grl�@^�!�[�i_�1NE���ȶ��ğ��������h�%D}Ղ �������W^<mq�ʭ��� ���o�l$���9�`e�ʐϿa��X�-�8X�B�2��jǏ�N��=�>_�,��w�p5�;�3��QL|�
�[��6p+H_%��W�3� o�eD���w.�W��i=����a7|/>�ﳢ�if%�T���>n��p���Og�dGa�ck���O2�u܋��c�{���u��r3�L�8��:M�s��}�� ���'�đ蹃B����)=t�l��:-��4�t�8B$���+����84�y�٥���dO��̰\�KU���ݐTY���Q]
_�b�[�z/�`(���,6�[rR~yz
�>�a�Q���>{�����p<����U��3��˺�7�x���J����8|�)�N��
T|�R��A����t�"�~�3<�Z���l7�y�m>�԰8JvY��L9�g�-F=n�� ��������j)\{M�}��ְJ:o��v ��#�nԶ�� �a��C]�w�'?��Pzc	v$����^$`1�_/OO�B��p��_��n�zt�����+��v�l�ռ��6r獃�%����	�f�Q���4���T̪�J��I��Rc(U�떳�E�&����W�:G|�ַV� 9w@� $`b`;Snd}���8C<<�R3/Q���G���yzi,մ$�#ݩ��QLbÄ ��" *R������娥3���s��z3���E_uG�d�=^��[�S��$���bj�w��4�Ǌ4Bӯ����Ǹ`�\^� ��5������.�a_ܲrܕeqv�z(�;���% �9B>H��l��(MWy&x>��W�tU�8=�^z�}h��h�
C@4s�_r���UD"O�1����أc���F�0(!�(c�QxE��3*l�̩)�0��t�H��Ɨ�e��MW����q!1M.�X{�ÍkM�Է�!�sI�K��QP����Sd�앶���V~��J����-����?��R��<NRȗ�5��]mK+�Nb� q���GH��F*�<�;�����e�Y��p%�1�w*�!�!�Ͽ>H$P2N��*D\|�Ƙ�懪��HCUW�z���A4˵o��U���w��Y�F���":o��Id��z�.k�2AL���6 ��y�_�Q�Z%1m����:��%����æ���f�Lc:$����e��|'[V!�ZЯ��¥���Ql=`4�-�v��F6��D��-|l�����T�LT%t��b��*b��=z��z���S�H��b��03��.�d�P�ȽΦ
���h� �j-��W�J�����|�:���� �P�$28�Fʋ��_J���Y��	�:NM(�^��+��z��P[)���d\�v*0��ܔ:��f�=�wIc����9�m:�܄'�|ŨtQޥ5�A��e����.�j� �F��u��FX�|x��e/��%NQ�xv�mэ6u�^�ԇ�H�v���!��2�"d*���(ZW���G37��Gݙ�/�� ?�lRXM:�p*e�\�;#M�SiH�� ��α�:�(�B�99B�l��6��{*谊�ţw�Oe�Q.�̿�*�v��ge>��+�#.UP�9d*�]������`IT�w E����ḿ�C�)����0)me	�_�H*`C�+�J_O�� ߰Z����]%�;ϰ"�n`S8n��u9�2�%��T���qdr���oy9�R`��A9�j����I���_"aU55�rdNn����*:�"��5�u�z/2��Z���a�[���-+R6�U�+�/6�2�$�ߋQ�R��Lj�X�+]��_������zN�5� �w�,�Ƹ���!/!�+2:h���Gqi���1�A>���q>߫,!� 9`���Rm[�
�&⍞�["k��t0��)w�R�MN�"Pr�Yb�@��(^�
F=��mΗٹn���bΫ�]��ތ���K�Z�ބ[UF��)����B���<��=#A�g�iYE��'q~�#|K݇�A�0ro7�c�!��uA�C�����$����z�e�:�ȳ0pVoV�T�%*�Scf��2�r���R��8�� d��;�|�8�pl�t{��И��W�R�41l������7�.}��E��e8��Kݧ]�~9�'��s�1Q}���4F`�l�2:��}�A,���S�*\?�S�r��E��L+��}8HkJ����-55��5����)ݲ,�)B���<�z�@�5/��K
��0?�w���Ѓ ({af/f��2���������<�y�,cI�<��!b�#��)D^�j8A���CG�g�"�[6}��h������"���)$��k�6ӽ}�i������4q������?n�;J�XJ�ޥnҙsP�h�cwY�AP>����-�|�_m�mCR����܌�s��7z(-߂8�ͤ�~�M�|}�â��A��o'&���	����nNI�����}�"P�#5 �n�������rA�J��pNS� 7ߔ�_aռ��[ ���'&tB'}�������x�\��L���aIЫ���a��׃dv�܌4�
�f��N�9Dѐ�|��(����V�|�o�=�MT��σ��l��mh�Q=�|B�;�b$��>Sb��m�ϯP6��>�.��j��}[Xidz�']t�=k��3����o�Z�M.��S�\��[Sk.�}���!X�Ъ�������x��A����C�si'����MXY

D�L��#�݅�&����"��I��B'�]j=�uE��aaA�z��S�$���&Y. z�� qM�f�M鸱�'���n]�7d|g�!z��:��"MOo��������@^Hf��f���I[Ap�-ԟi�x���՛?+	l1�tg�$?N�)D/��d�0Cj{@ ��F��Y��>��(�\�\m*�)�6�ex�������}!$Rȣ��c�ۜ�2�uӯ�A}�e�oN�&���_x�Ԋ�uc��Q�бy;o3�؇��߅��$�h�s�W�Y���'T��qQ��pfS(7�';����Ӥb�Kʟ�9�dqE>C�9����̢Q�^�ub��"�jy��j����h�f��6$νV�b�4K�sSt/_�q�t�Dy|�X�X�	��k�!Ƣ�L�P����Y7~y�p��Ez�y�2�r\��"��!�L��q���ō2��.�x��Bxq� ���?�H�{�*�`���@b���ac�2P���^�B9X�E�m�\�;�^M	�;�T���9�b3B�1hW3���g��7�V�����\�R����A��k�'4���؅P�F�����JX�.@_�X@�om���9���F(@Y���k�t6��u[�� yG�f?w�X�ko�2�+6��9�*w�qQ�N`HQY���T��vsg|gJ3��o�|���/�� ����{=�!�v٩����)4�E(������c��
ٝ����w�������jd���w���T�g�>���;n�����]T���Ae��[�=��C���n�N�j���"�� u�-���6}x�Rv���<��Ѳ�Ϝ�Bm{��xP�m;.��G}(�G�L�
+g{��\����Z�B�=��%��
yXєt��T���[�K�˩���6�2;V��.��B3�^�;Lvߘě�8t ~�>�	BŹ�։ۓ���ŷXF��^�*R��۔Yp�+Y��,����#�s�
;A�>m��@�E�c�ŝ�q��I����
u��8������֢|�r��D��Y�j���Ź��U����p�A�/�G���:����"��P&o�!��P�eeP-��N�9��dS�C*��<ba�͚_Hi�{<@[�wB��<uLn[pPxٸd��9��#@��|M,F`}d�e;w�F�7�{(8�f�QI�!���И�,��_�7�n�l�M3t����1'�d�4�Cze���g�a��WdJ@�}�����w��d ��go�տǑшJ��@�s����@�������Φ�^��W�4kv	�������Ad	�����"�4	����}R��?ix	b�P��o/�l���t)�G��xn��w,��g��U��."���'i34�̓>���)G��O�]V9Tn���WVm8尅Z�j�Ē���O<5��o0��H&Ea+.��,x�
�x��#�W�Ì�Tt�y';B�]�p��5E�p�C�'����A(~��QV�b�f�n��$�7m3���y6CD��s]u�"��PY,�B� <N�̘�2�>�-v#^�ڿ6�)�g-�zQ�~���DF�o��b'۵|��>��؂�'d�/rbE�r��2�T����r1
����&���f;MZ
6��Q|���b-ȵ��������b�8��n�ۂ�c3>��mp��ãʽjq/�)x�V*���RG�-~�f]�L3>�I[���������R��"Z����:ϗ����0�T�U�Z�C��nݻT�3v�q<����x��馭�^"���S�0H���gS�v���
�u�!n�e��u\�������M�!h�s�\|�������`��oOQ�z/j�(�Қl��Üd�1�Tǡ&BuC
�Ț���\a(�Z3 ��_�
�
��f�r�?k���ǀ�ߐ��A��刧,"*����c>���zFfQ�K;�OO)80��\�F�y�n�}G�Z�%\�hÒ�]�j��^����qː	�aO_���T4���Y�R3d�D��U�	s���K��*�@=o=_æ#������!����)]i���` n8ğ��d�z��ټ^C��#�{����T ��u�/k��W �s\���@]�v$��z�H�x�վ������u]��+
�A�!?��$����E�J�0ͳ�I�R�s[�V7�hJ����Fi}���'���_J��a�{l�ȥ��;Q(z�IV��XԍB�L�s-���.u��]w�׀1���J�����v',#�������pל:�>�m�6^�VQ�8Fz7EmG��Vޢ�܏\ϣ���<g�\.�����n���d?,�ϟ$���pإ[,�(�{�lUJ B>��uK1?b��ң]"�_��|4 !ݲ��c��r��Oߣ��V�!.���s��w���>ZDٱ����z�������C��!�6�I`{d���'(��g��������6��ڔ���w���KD�r����+�*PK���;c��>k���d 9�����Z#�/U����ٻ7�8[�9��U�|E�@m6���L���Ө<.5���"q�/���+ԣ�}��X���Pg�۵m��~ӻ�d�3z]$�Mxe-S�� ��=��7hv��@�$�G�<v�Fq��:>���v$�b�j0����̜�����5��)=��:�-ʀ����ど~���S+���Ȧ	�5Be<;����"����9:l�M%֑�q�kX��'��O	�j����e���7��F�68�Ϙ����M�I���0&�eؗ�4�,f������X:�����QC�LU�x&|�Jq�(�r}L�F����Hu��>s
Ƨ��cC�_�v�K��������DM��1�$�ى�]�Z��2�h�lmt��b��?n��o���h�n�IW���r`<��C�V�X����d��O�I�P2Օ�AQ?�rj��RJ?9L��J.	̩K�&Ad��Jt/��5�|(����*�6�ipZ�����P�'2�s�ބ����s��Č~�2�n�d���v��`"���+���x|u#���o/�4v�Н�w+�ї��p�����Nc2z4�U.�J�T�q�_Xԃ�Ģ6��}|�5[|��R���.��va2	P*t�{�@�cX��N�Z�m���ў�0���:�쏞��M"�_�����s�͚�S��k�y���rn�ﱒ=���8ֳ��,�a����q��sç�J�ZY�?��P�b�Mk���D�G��|���r�h��X�
dMc$��^��r�>�(X���REN+��*C��:3w'�f��)�C(�T�E	ON��|�]�]�/��aX��,2��C�beJ���Q��Ǯ��4������	ˣ����5	�L����R�lF�LU_0Y8,�7�����.�TH2/;Y�����t sߙ�e��nk}ݫ�J���&F�E����Z]KE��df�InPA�7�e[���� M���D�@Ҿ�L���9�f�������G����b��&tt:�6��"����6����= {�N^��!�1�??�R����)p��']Nu�<�\����b���<#�|�)��+��%�/�R.�fJ0z�@��i�.�������c���� �P��V�C�~W�5����ח��U��8�K*���a s5��25���1K\A�Y5L5�����d�~5��{;Rq�+��*��S!]�GF�|I^F�������!�$���mؾ���?�1����0��ш����Ȍ�Ǔ���>����BнŁXc+1�����2@<�� 2��̼��Q����1*}K�䣽�/����sA݋J���nl�Aw��}|��t	�ș�Yo�K~N���%߻�%��K߰�4j�ɧ}KW��yN�ԍ�la�oP�����2�X�<A��vE�h�����{d���K#_��$m<۲�6{��(C�3����ƅ����)��vZ����)'�Icg������/!����r���:d�+��`���e�, ��^s��zM�5S�T�g��$�w�����婮�;�쫜�iΪZ�Cs�����%�S��r�{V/�-S@���~���P5WRr7Mi��H����:"�0��MB n�u
���	�z����*&]�{�3j���~Oʗ\��޵_�)��A�z^�R�` ��Ïq�(��f�s����ФP�vC�B<�(���N�C������l��gb^�}
YR�Y���P���&1Uy��մ��C����oX� �i�v�ɮ�����T��,lB�׵}7����5:���b�B�ζIC� ��rL�TA�v�,���V%?�'�Yy_�|jBd�+ޒ�@>3�7g�V����rAS�roR��=˨5�,هhK�Dł^0k���`�x�,��v��[y���ָ�Fwpn�u��@���g�6.��OIV�؈�b�}�2>ݦ0�=r�iL8T'��[��_���xG,��e����8ُ���Y�һ�&dx��B��md>ͩ3�i��eb"��.�\��wh�wR����d��ԩAF�ኼ)��r���bƮ�H���XB���~����39��C�r{V�2۵���X]:�޵���&=�Bxk؈D�F��3Pu8��k£���{1�&.|º�1�-H�o6���������J5��� =֡4K��B��Y�Z��zl��Z}\�B���>�/��,�!NAn�Gd;C�;��[�����)A�UY���n��#�d�����^�Ҋ$j�F<^�	��E���|�D��j$��&Z�	g}v1P��;��4,�_�b�-���T���v�(�Ky&+���v�e���ڗ}G�B���2ZQ�|����v�K��~y���I�,pM��d�ϞA�te;��ى�Q��b�zh�Vկ��1rdP�����Y�E��m�K�)w {����zğ�-�^�{��rS��KHPGU������N%�����v ���9��δz�P҅���� (��oM�;��U 
� }#���j���_���C��ys:��Z�������2{���F�p�ێЅ���L��
��!����&'Q��۫�����*�D:'��_��"���>]-���"�'i��b>�[4�cЖ��>d��&�/�<�!c�1���%o;C����K�I;v5�X�5d@��T��i
C�նl|+ s�n��'
;��[5c�ɍ�^����(G����WFo�V�֣qۅ��cyG6���0^���
2��j������Bs�]W�Qoǌ���2�b�@�N����>����o���q�c�O±bᙔ����Ʒ�����F ����_Zzl2��$�迬���#��o"�W�ܢ3S��1�|L���"Xj�c�m��.��A�A`�H����F
�ր ��w����|�^x@H�E��ni-9�>}���,RF��[���|�Q0%�-w-]2��Ai}*hݙ�Ef=�L�^.3�˃�P.qE�,��$|)�!�幩Yj��*�>����V��9��aZ�3����&	�ŷR���cb���$g�6��l4�I��'f��h�:]�8���z1X���ǃ���QAM�`�ڈ���6u��3�ò��z�U���ZxOߞ�HR�:ҙz��T��1�)�����z��J�YʯY���w4%�C2�{O̿�Ah��D+��'\�+�IT5`0'�//����ڄ��U&�s8�/B��P8�b�,��&��"Nڄp-�����@�Ψ{jY�to�ƿ۔�Q�<�`R���ʼ/ݘ�I��)�li� ~�g���4��^-��F��g���<�w4��J�!,-6�m��#$3Ьa��o�kO�������R�Sb�H�06 ���A)�d&-��P,$�2��^��Q[�7��#�LH��i�/�q.���\UxW��t����PC��/Ы����饹�MF����ʕ�j�����1o�����_ލ=���o@��H���I"W����'H���;� ��� �|�Gw�Mwל0%q������ӿ�d�ր�}�'�J6.(�	�Sۑ�\�"��B�Pkg�U���)�Y� �B��b)���E��4��p�8�>~=��8�Ҫ£��
$R<$ /(�'G��ޘZ�[���hD�Qaɽ���E�aN��+��
U�]6����Rmx&P� _��L͏��� �������J$XL(����������S�s�[�al�	��F���I��W�`���@lK�)�!�q1�4�|��*��2� ��}r�w&I�G��V$�ݑԽmsY��8s���kZc%�$��I�?JN����_q��1�>zzq�����C�E��x;�K�o������r�>1����`
�-��T�΁}����Bk�	�P���5�8w�s��b���T������+�}j3�Y�������\�{���<����i�H�����e̗|,�Y��,�ی�f�W@�|�b@	dBnZ�-Y֩W�֦���XG�Ī�A�8�y�T�T=��'Fѝ��0��u���u���y��h�В�c�Ӟ�&R�������D�n9((���Pb���8�҇���D��w�7-%w�F�(c.�_���[�ߕ�����z��/G�日��7tQ#�����'�`YT������Q�g��1E��+rg��.�Pm�ʇ`�{�r`]�q��S�����T>]�6�~�$#w���R����	�m���}nۙ�5.�c����^�G��e����{���3��Ĵ?�e�S���Ϊg����� �q k_|�C��z@�9Z����ѷ㷵wK����득�A8����!s&7�|o�w�����c�;a��ʕ!>_��^��i;�H�R6�Ə�]�i#P}���s	���{5�����f�Q=q6F�$ujw��L���dx0����y�m�*�*zo��,�V#�)?�ɵB0A�1�fDa�Ҹ����PD���������z>z�l�r��;�%�!.:f6z��3�$T'����{S<i}�	��
.��5%ٍ��|�q��|�"��ʉz>�(�l�$�����u��si��n��Fѩ��$ �#O�ش�HLK �n���:,0T�b&jk�C�]�Z��To"�Zag��I��AW��{-`�Ne7,t�3���G4@'*v���2��C��0���2[�Գ�ي��M%P4T���!�Ӑ�t�+�M��@t��A�;Q����}��E �V1����86��h�W��@n��^
R��n &M��A��ǐ{�#�-b���7+�4���@>�\��G:bZ��Q�^g��h�f)���mw�hP_Nos1��3mw�Q��Z�a3���7>W+�Aq{
���Q�|���J?*�2a�T�:�fO�W�LFۦpW���p�������F�vb/�Vؕ�5�>E].FZ�V;�}z��Ż�	^���"��i-���L��p�i�sCE��^���U	2��<DX��w��m����9��'�����q�Gjk���}O�����`'�Q�� �!ĺ<?+1���.��4�7vjUĭ�Ԅ�� ۠�\�T��	��"U�<o��z���'F�f!+�	N>���ת��#��ۄk�EH}��	��3�����_6c�K�������Pfv���rt���teYmu7G��[hPsl,�5�Y&ڔO/��7#����bŒS�!��#V�\8!C�/#�b'�<ޜ�%ԉ���%�&wDp�J�3$��
"v�y��~��:�D�7'}�a��	E�v<��^2J���S������د|X@G�>I��o��E�c�j�$�`�оY�]
9�5lU��i��JR����jFN&�"�3�DyW�^�?��Ok	��W(Y1�ԟ�bL�F��~��|<�"�5r5}?� ?��q���� �����M���߶�A�O��:�z���J�T���H���K�q�x�I/��y�I��Ą�W|Xxt�����q裓���
BL��(�K�����{3�U�]!��k֒'���Iײ,YSR�c�}�w��(V��0���iS!���Vb��^�%y�({<q�X�RC�sk�!+�UM�+�C����m�K����&
��ա�-`��>� 8�Z_�<�����y`<�_؆���me.^�G���A�X�̈+����y�5ge�k���9�&[Z(��p�Y���Y��E'#Ԧ���Ʈs���$�g�sl%��e�T#l$���6X!�&�5Fq2mm<%<���{�P�X�1�,�'$ɺ�Y<�C�W`�82ur� ��WnJr�m�k���e{�RZAi��!4��s���E^[�x̯��v��K�L��7/u7��Ri�7u�t�������������b�k���Ec�ԝ�P���f��##0�`����"7�9�J�s*��fXG�>��3���s�ܭa�d9�	J�V&���|�j'&��>sk6��p�ױ����.�w��̛ҞJR�N���4^�4�"1TV0"ݞm>�6Kn�tL�)�V����i����Dٚ���Z�%�=�8�Yz-"#����d�۝z�]�+P�T��t}���gX#��flݓ1�n��ȇ�a�bG`^�dNL�MB��m+��W��ߗ��S�2�/���wX4(
O��h�	&��z^�~X(�ե,^��~�'8v���o���g��i��7�d���/�ȐF?ؘ/��l��̬-h. �X�&-@��-��z�5�-]N}M����l�Щ���n�fժr}TCN4�y������K1�v��I�*i�4"�996(P+��BZ�#*��U*��z)��'S��2�1��)�1���oQ��?��F�e�a-�X�?Vɚ�躀��k8#�]��y�����pf7�����P�͕��B����=���}��Zmj���χ3� l;����,O��ջ�K�=���y2�î��s�z���s��������	mr��KHM�G�C!�| ���Ζ)q�d򋑣Nb&�c��kPjǟ&�S��Z��I�:"WB�A�S��#ݹ��[`�pqJ��
�=�V4����YqB �Q�e�N����^�� B���K-!�+��BQM|�	QY��hBvT���_Ԉ��*2�TRg�D;���r�R9�7<5�u�3���>e,_+�Dn[������18�+CP���iN��Cˤ�u�٭�Q[���s���u9׉���WC9��F����YW9�ps��vyu�˓fl��9OlU@17?�_T��&�z��yzf�p#��J��d�����y|�Id�.��$"W���N�Bݱ!�Iv�JM�����׎#Y�_M\F4U\@c�:�إ�ul!��I��һq.P`��Tn��ԴSU\�m�%I���~�";5GJ0�|�*�- Lv*R	zѿX��F�F��R�>�XF���:�n;C�al))ҟrR.�����!�y<�a�ʗi��'Uz)�hp4&w�Yt&����d��|�d��j�@h2q��9��xJ�C�ՔO�㝄��"~�!2�5ǵ���~��cWN�K!)��1aq��I塢��^���eƗ�76��)�z�L'��������ݴ��q[����� �=�O�"��^7������L�pJ�x5�R�բU���X�>��7�3��:�c�deʾJB��XI-/ns}��\�0��*V�7<ـy%ݣL��o��t��󴮙ϸ	z��:�ՅҙU���FJ��0��1&�n���>����Z��∉½d����#�h��	�y5���\�D�C'}ހ��+�6L��X�����}%� ����������W�Pd��_��o_+D���a�S��o�Q���Ӊ��4>b��ͭnz[�C�G����/|���)��e�~�L��Z�2b���� Atigz����HF�\r z�XP��%�%r�DT�f�����/ G'�,����Zc�t�I��BWfG��~pS��k0����[I7��Q˽Hl�^.��9��X:��BQ4|�����#4g	j�^{�ə��6*�*mR\eͪw�#�*�@2v9���$"�߯�<.`�V�S�d��º6Uf�v"�t擸�����������H/-y��yܩ%�zz�!r�%��)�����h�l�y�]Z���Gm�I�V1'�}��rƃ���TH���Kz�B%�:E-+*Ss+j��/lDq�Udi(5<�`�Il��}1�
X[�V4�ڞS�][�z�&���A��ǚ$y�&���V-/��A�}	zD���u�����t��"�j�e�N�+��DR���Q�rv����ƶɧ�(-K��L�=��F)r_��&#;[&DS�#3�f6Fш�Q'�Z���nyw���H���G"�C���m�4�+�(/��Û�8tge���`nP9
Ε�K����<}�J�(ϵ)/G[++�9����@�k�n��fAӳu�BY�d�s�#ȁ�^�|���� i㶹�z��
�$�}���B�����ƙŒqz`��x��a[�!A~9SQ��Q9�W�	��>�2y^���n�g?R��� <:q�(��?�Y����J���H\)�R}����᧏�禪��*����v�&�J�３�pςwT�u��ux=����<V���f��_L��w�Ấ�
��<^�_��a�g#F5 >Ӯ#�L�@x2��ˍ��1�sLV�#��w��TY�B��,碯�z���{F18��*ob���x*g���a}%U +=_i��U�+�?u/��p�g� hD��8�V��Ít(�i�!)��|f�c=�HI��6ô�G\Zi��y��~j��Y:=���1o\�ЊC<t�CG�bC"wd�O����6�gpMF8��|����s>��_���}u�o���J����S�O�����_xy���>J�;�����U���m��X�m���Z~f��`M���J77�Uo�b�a�����,� �[b����-��A{�z�BՍ��$Td��O�E۹����k�Sg��C�\�^�	f;eY�$���u|-����o�]/�!�ڦ��u��㮫��@�<�����0����h�����!#�g�1�;�gZ t	�+�Zp�C�(�($�t�*9��φ�(�܃nrSVŎ���h�V@"��kq9�����W�(�#;�o-�<�Z���(�s��̣oE
��7";b	��V�4pJN~�J�}avv,&�0z�sxR�<CI]{�uH�S-Y݃�T[�������)��'��#�`�����\�l���
��c��R�^�W����L��a9X���QL9 ����kU�ql�|C�^$@�&m��7Gbr�M���WG��$IqDޭ�2%}�y�Ƌ�#�R�5�t@K�xL�h��=�O�8=x$.��^�
h�����2��a�h����2+����yHV��
4xJ�$�d��H	��e�w*�D�Zef�I�,��W�Z֍_7�|��.��	|�EШ�
�$�����Nk3͊U��Xj%|}����?�]܌����E@�m����پ�+VcwP��3����w�V��@Ef1ؽ�h�k�C�1��)�;�W�|U^$�qMi��+�4�t��+��^u�w������������jge���m'"��D��|��ǌ�4�O�o}{!s�93��Y8*�t�k͔�9Zv�QޮR�}�x�<��c��
���D�2�Q�t`��a��"�+ǆ���%A�&����ʼ�/����֔ҋ�y�R�L*4�^�\E�k��!;*���U�.��*�eN�e�5�2f�r��n V���O�'1{u�f������	4w�1"2)M����P��J�>vn����T��\߾6U.B�_��nco2�� \��H2�����dI�"kmrm*,L�f� ������fȾ@��g۸Lny��_�ΐ�`��n�#t����anVKE��"6��﹆+����T$�8�iƫ��@c�0w ���`cГ"ۨ6�]�*�w�w���7�́�GB�^&c�i�91������(L8|�6Թ�;θ!��`Z��.�y�J��(����.ۼ�Ň���H#R�}�����S	��<T�x;Pc�����"H|N�Po�.�>��`�}Y%;������/����aD����%��I�C�nE?�R��F#Su��������h��C�'��������:L:f	Y�q���TK�LQc�i~Րt'p�}�r�R�ۇ�C��;Մ�J�rz��	�=�.D�ac��[&i$���"/5�.X��j.�˧�iB1
�2HB��Rg��Kϋ�f>��:���6�����O�6Ըs�]��
�B|�Ǘ�C���� n!Sۣ��L�}��&���)ll������{}�6�cюPa��h�[�5�5Z����՛��"�I��`)o��Z�����V�bH�G��#�R�G�s,9y91�)#�y{Z����'��*\@y�q5r�꾚��yt�zK(�Ȭ�2�0	�� �X��4k�gat���������A�"��r'5�~��Գ��.%�m'M�Q�{�#���G���65z�,3�����G�J�c����J�Ph,���=x�I��X�1N���1f�qL�������z�^1�r]$S�:��z�[���� M�Zb�N�-	�k)�����
 ��xF���[J���Y�%Az"Y3�*��{Cl��(0��X�_X�Ʈ@z�ܓ����[��.���	�Nt��5ʊf�����rkc��K�ɽ�pj����@E�&!u�mk<S����-6����������uP�~�1&�g($H�(-��j���=�K��Wþ��v�$,�U�a�l
�s#���o�6��4#��S���}O�V��_H��R�&�OFs!ؓ%H�vZ&s)y!�;������; ��K������x���k��nb7��dW�C�����T�h?�f<aŢ�;��,�"�@�h�Ҷ���L�np���z����^��^ʫB�%��@��_F�e\�̾O���~@�Y�.,٧��,ג*-��9xb4�-��*�����љǟe�d������s_�⸇>.I،��:]���d���0�����,щ��	����*��6��A��5V���:8�G7�	�����3��l@~|bv^T�>��%�x���1��(�������H��2�����Д�W�}�Ez�k����ELV߹�ݎ,P�Er��¡��c0b�BP���v�rIư|0���~XF���U`�����Xޘƞ����1�G4��_�0�<���F+B����u��G�GӬJV�@pqX֡�m3��Oʖ7Pl�W��c�23�/SU�<Y��i$��=[���%�+xa����g�J�	B���Rw_�"L�33�w�L����Ub��L��S��*x�W�w��ɿ��]Y�ֳpa1�P����#u4��B�����S'�m?�ˀ�y�V?g���8�مީW]�$�"�s~Qx<{�?�P�esϨ��U���ͬ�򁯌�Ɂ�q� d����������5N=�2@5��0ե��KO-��Q&�����ry�B`D�֦���'��a�Or5�b��f�ŞyT*+��Xe����- �s�:5�� 麼��P��f�W�j��`~�S��ru^L�$��-�d1���h`���Ň���	�X�[%8�J+�Gw�Euo0���~1�k�}%�/Hz����T����՛Q�}�m�;��:޿�8��}V���
��lU�5�<& �'��Mrh��b�$?�-�+ⅼ�]A�3D�@>̷g0�=��O1�m �e䁊�^.�L��aW�V����� ���K��P�!Ĩ��TV��G������g�cޭ���Ǳ5�1u?�-���P��ŋ�B�т�ᷨi7�ȘQQ*4f � xG���L�����D�6 �}>��3�/�r�ժ�D��}!�q����Z�8j�\o鎙ȯ8S�b��B��~��AF�uj�W�k��Kz?�)�Vd����Pkf�~����Z��iwٵ���'����hp!/����%�L�r��eG/�I�̖3�����-��P'H��"����S�#}[$��Ll;4�Cǲ�I�G}r��L�JY�up'� � ���{VGህ������f��~��������1 H�8r�(z��Y��~��.���"�F�"'8'�"�joY��TYn}�A�t픘"��c�}{R����5�r��O��g�4d,E�X��Җ���i '���υ�, ;��.8�U�${���e�M��VrH�7i��r��g��w��k:�R)��|O�gl�u,e�<i ��3�U_B;?Mj�vˀI�8�,[�%�"wSF*����]�9��c���+�[�*B��{|�[:ݱ/�i���9S:>ѩ�������9CW��"�+s�Hd�t�V��o0x��tM�`߭"�+����I��@�|���^>�����:}��r�����y��X;�d�)z�)D��[������α�|�ԧ��N
Wx �$qȐ�ذ�_�dbAp�.�Jݢk�#�Z���f v,p���r���V�ş����:m���L�_	D@��|�bw�`Po�.<6Nַ�[�6'�m4@]�l�㴄�E�Ko�ŪtT���59�𞤝��Ñf�9[ӚB`�q?�ZVg�G֯�a�����<YkMG^��P���b|W|>W�VQի��{i���vN�%܆fZE�+�H	�4%p}'PK�w��]�y���`!v\9	�o,q�`S�:ˬ/M;H����SC���Y���m6�Ɵ�a��!w�J�B+eҹ���Inܽ���c�%2�C}Q���ɭ�B��V�q���qv�A�+�s�+g^]�4�|E�Z�.؋J��Y��%pV>�`���:����SmH���0�������Ǭ�P�j���6 eNH����_t��]�FE�8��V��L_�i,a�����4�u���׈GCz5����jK{�h�}��.��(uv�v�l���t�i�	"���f?��x�j�HΔ]�������9���@,��0���ԥa^����m/F-�);�=���~�9���7뚴&�;(E��Ξp�.Ъ���~���������a����>��X�m�����
8$���J>���������	  �$$�c~�o��x��y*�#���{�WB�S�I�@4;<���|j�1
�`;ю ��"��
+
+��" zWx�i���۬�F9�CE��QD���NB�����w�o"T}�ʎv�#��e`���,� t)>r�u�Z���s�����œ-����^.�Ay��.3F�-�WT���'�⛟��J�R��o���N���1���L�	 Zi"��<��(��S��؊E�E*&2>ۃ��o��Z�� B�b�z���f�d9]w�t�G���Pm�̗���YU YP��=���j�mb"_��C�<�G�i�!�uҊ��[���Q�� �6ӝRJ�+{i�����V�>f�����]Ek��Ѵ\��k��1\]��qS�ɇ�s�p Rl����c�=+�衳���z^�`���2�cy�K����3����ԙ�euu�;�����h��%�Ч���A�D����!;|x�n�i޴��0H��=c�[��s�p�����ꔪ�uOI�f8�GA����5�O���8Wȃ���	�z�	緅O��XƔf�B��� ��gO>�M��{5YI���ByDU�[�/��t�����FF׸�}�l%v�ߓ��(���R��R���>�c���"� Ws_�e�(u�~�u���ⱓ�}l���rO���sb��/2f@�`��4?}�Py{;l�~�ѽg�g2I*��\��
���`�û ڭ������Qi��B*8����t�|��<�,�24!�7�[����@h��=~���'4v.Pi�,�'�z�ѕ���tr��]G{-x��4��6�
e艓���4�6M�JW��w�S��"�$�A]�E�}�0�$E�J���=�j�cN�&���:���g��u&�2��.�*#Ӑ�Au7��S�k	�-�����У�Xv�ў=�L�&�����y�h��*�o�@���<k�~������h�S�����ngS�O��Y��ԘK:��]�XP��7�0��V�1 �2���5͠Ow�ob!�D�a_�fH
���C#��2�l�ft�%�ڿl��p���ԓ���·�K��jr�fp�ˊỶ�!�9��aߎ�:ϗR"W=�B:��T�4�A��l���ײ{��Wô�-�3d�S�!S�
h��F2p1��� �_��'�	usH��B��#ٮX��D�	�J��@^ �f�@$�-f�ؕ{J:�qZ;o$�cMVk�7*fN��fO���T��C�UM����}�_�7	�8!u���3��tx�ৼl}�}�<�ȯ�M'B�	!�^�(���Y'��0q:g�!�D�q9���;G���f����V���d��e�:�B{I`���M���`[��K�<u��p����o���kH��H����
�����蜀L�ʘ;ts�D~J
y�����F�`X#��+�vx}�qt���fs��S͞\�$�CP��0���x5��>j�s#�l~�I�{�H���~�t��G���o�I��?-�Oh�Ӹ>Q�R��M~�`'U�\k�W9����e_E��JA|s	���qŴ�W&����I��B�%��r���Fs˝�l���[�:��9��_ʸ
�2���5@&��\����m$ч�aO�=#��U���f�q��MeP~E�ebF��}cމ�i����	�9��?�j^��2�r}_:��&��2e�¶��&��)\ CA1˓�:�f��[l� ,�+�����醼|/��8����`��k#嬆���ƑKM��,�&ׅOL��R;���x�N9Q�~ьF�T�dJ�� n���(,ZV�K���^�R�N�':�,���eiU���A��HҟN�L�'ٜ�V䬛x<�!��!�]6��@qZ�s����H��G7� �@J�E)�F��	�<�=�|z�+��@��T�Yd�*���a5oD保�0��������N��E��%��C�791y��.Tb��N��=��4�$�n@r�;P�,k׺N֤l�m�:����W���ڼ�+Ȝ���D�&�ㄡ�x��BzϺ��k��9�O�&�<��!7D��HA��T|i��.�Fe r���+���M��W�mx26��g�g�>�O�H~����ê�u���
^t�
�ѺT�Z�O�e0e����?�u*��T8�.��*qg�[H/KQ��6�M������*�;.�sZ@�'*7���dx�h� �ʹ��g5�\�fG�$���u�p���8����_
05�]�+Tb��R�w-'fbBͅ�Y�*��۶r�B���q��V��ꔗD�\�I�N��H�yC���7����ʄ��&KT�C�~$%�<(�� 2��z90��b�$&�i�6�f�4�\@�a��DK���.�/&�@��h4���.SY��3��>��IC��C�L������������{��o�p7��2TlU�R�?�F��%�)��[��}��K�Q3�<X9���Wj�CϏ���s!&:D�U:-Vދ��+x��&z������f1>b�������x#U_u�� f/�92S��T.�4R��M@��섭����~N�)^�(�e�2Ď�(;�;�Ԧ��Y��0j5�z)�N��Rk��~n�S9�0�� 4�p,�����o�lĠ����
߱٦�^��@=N������������eh|u��ާ�о��_*�YM�q )�LK�ʢ��Yk�(��G��dO��7,�/5N����Q���&hԔ2<�9��������ǫK.(�����^�"]�X�Ϲ���u�e�O|w���s��@C�W����g�GQ��7]9#����g���`t_������7R�>�&�I���sC�c�g�؇'"��Ͳp�$[)Lؚ���VT��є���1@C�eD����o��ڵ���i�C|����8PMxo��9,���0K��f�n��W�ߪG�$h�:ݘ�L�����������BĪ����#I9��'[�%�k�n�pT4�
ܘ�u�Y�#�.��f�z�?ˊ�!]p�tu��x���%�x.��T���ר��$���rz�B�~d �2T��q/��<��,�q���«��g�U[.ޥ2���R�u;��1�&)7�&�p��\�cx'm���1�ˍ<bx2�`��\�Q�"�.���IyJ��.ö��<���I�T\`.���U&�s��/-k��u=Lx��jʸ��	xK�i��PЖ�>U!Ռ��u���L����k�.��ߍcw�ҤC{��ɯ4pvհD�C2��_����+ƫ+U2���:N7l��]���vl	W%����V[�U�*��8��~��ר-q[\	X,��Nx\z $l���B��fW�����L  So�|`V_Χز"�5�����7�0���4p"�cKKL�P���I��|q	P��� ��HI��o��s�$8N���@0j�M��ك�*u�~�Ӥi�?»�Q4�-�Ό+�_�UZ�ˁc����,Q���s� �̆�i��>���s�~�:�����&F�;뷥��5��������ɆuB1��됂�
r0F���J�?����@�I����aa���Zц�J�-E���̙�1�i���HŻ��k-���+<}����*��@m�b��g�&�R�0I,��S("BV`nd����z��v�u�k�����\���Jc���J�#{�)�e3�e3?�5L��B�=���}y��`���5?%R
T%,��O��E'���hѽJ��z�����~e|j����2ִq�:��Q���F1]|����=��FJ��F�{M������ƅ�߿��ljo�]�6<$/�=�|-�E�4�ъFM�Ɣ��������k�HkנWe�/�q��CL}}��`���]��n��|i�)��<�gd��(y�1=椳����n,���?W��r�3��=��]E@��,���x��S����5���:Ku��CJ�
�Nj�>��D�ӱt�������X_љ
�ւN�?���yR�(���1Bgs`�r��RF
��b��X�Ҁ������*�g�����1�X�M����bA��yb�Ʌ�|��w毎>���9PSAnJ��S^�S=�Z���(��������v�`����&����b���S��@�%���qs�����R�# ����d�9��fP,R�Ĉ<��Hi�g{�XI2�����r:��{Ħa�����i>�+���Cd{�ښ�03�qg�CO��[D�r�<A��G���M&�,����!k�`4�C��\z*�����u� ������ڼ�������j�-Ӑ[Q�&�����.��"�ev�聰!�h�k�9�CUS�w�$2�6y��������>��2C���l���fZ
�|�e�Qc�%��R԰>FxLb���ef�k���1�Mm���z�����t��	xO��=?�����DK�0IM��2�����}�R�\<A_�1ћ�థ�̺��ʁ�#� QzZ�=$P�Av�4��	�w^�[4Q}#��kGS�����9�]�ʸ=���`����	0g��!E!Sڲ�$\������j�fWsˣ7�#���5O�ܜ�3ZE�I
p�T
�X\���ѹ7�*��z���SvO�_ͣ�1�:& b�j=,�[�åj��΃��L����X��4��_��q0��f�)*����A�ohuv��؎�7�/WU��F-���f:��ߩ�'�����`��+s�,r^
	K�DY��Q�D�¥�͎Ί%C�o
֚/�,��vя9-}��c��_&'�Ԫ�U�t�ECy��eg���
f��S?�͒d����)�jxj�sM�ydR�h�,X����u��T��VT��N�I,Q�s*���xM�{
~����<��sH�	�X�E5�0� ��2���2����CNJ�G�������%(J�� ��LJ�q�|��	Bʕ:�Y;��Lդ���Dǧ5�BaJ��������LOy*R�'�kV q�4�`c�4��|����T���t�t� �W�z�/��}�Ź?�����0D�O����������"{��][m^��kR���#��C�kdn^�\ߓ�>�#��_n�A������'B�xƻU>41k�y���E�4k��B��eH�E�
>O�SU-pC�V��r�W���$�N*��M�g&ښfJ?((�J0�����b��M�/�����;�,AY-,�_��VOV�l�D�v���4����;�-yEqB����fo1�����SU�L�+���`����1Cƭ�%�3g�yqpM ��1�f맟��c#`$�l��"Sa���R%��if'9�}��y��_�f���Βx���21�P��]Lk��*�?N��S��*��j�#�а�x~��6����A���a�r=H,>���Oͱ�bcsA߀j�$��0�vf�w��>�� �1J#L�s1<f?�E��p%m~o-�F���e:OB���١ʞX�s�T9�\�>t>��g]�]-�t�~�t�b>O�|��֚i�eW}�=o�9I��.�Y����g�_B�������>�G���{L��%ph?��ATBڕ,h�Ā���sЙ;����ӔyKr�ߵ��S+0Z2���7p����)h����ZԠҝ3�o�s'M���ԛ�.�r��fz��^�.C���D�4���MD��8���Yޞ��XFhܚ܊��;5�OM�De��lo?J��˄�����W���2ݨ����(��6V���!��:�'��1��9a�������}ź][�"��*����F�%}��.%����-0v���⟓jM���]*wJ{�i	����wmB�_IO��Mi��D����iIC_;�g��l��X�e��-�Yr�p����o�����$�	�_h/l��ђĶ5��@�!�镇
��*�e�<���P�k��3!P0����%�t���#�F�`�Fm�Q���n�R��]��d�5�e�S���?z���Д!+HV�FtK��hPn�b���s�b�a#��DK�3�j����h�&�cqE�sR�Q0�8��ƕ�~*�ލJ:3w��.�̓��@Q~��3e h�Eoo�8��YV���h]*�Tm1��)���[��T$�î^[n���z�|v��@�L�^a�ʟ�Qj'���V����h0����&pc��44x��s#=�4��A}��{x�d���Z%����׶d�B�w��Lu���@Ae:Y=�� sk���<I֒�K2(jt��k��(10�B�������@03ƻ������3љ���k2G��J���wvo�G��$:#�^����!^�E�6��3`�����+�!�2=C�&b�<���<�,�,�%dz��Kb]��.\2���B���ţ"��Ptޠ���M�X3'D��5��D��N�T�%)�;��`�Ә@~���E6>_����:�5��^l*�Z�#����W�aiu�Z���Q������?ijºV������:�����ɛ�2�9���������`�ӊf1j4�Io�c�h#��J�ak�Mv�W�`�A��s3�/��O����h$޼"�n�(�iֺWV'0�0�*�W6T>AHК���+Ie����X�Vv��7y���SR&�/�N�F�_����,l�~>_-GIW6���Z��J�i9����(��@n���,Q�;@Qq��Ko��m��*���P�_ɥ�!V��I�z�?�4Id:R��cU���:y�J3�������^%�Td�"q-�M�M�X���fz�|�}M�]_ɎJj����\�Нg�� ��8���E�z���C���
�Cg�`Qi�����d�����X5��[aP��lT��=ߣ+�~��F��N�a(\S��9G���?Zt��.l3"���h���^*,|)�F@����f@�o;fW
�i�vh�0!gt@���/)�t����K�`�n���($����*�%	B�m��̧(����iq�ekʘL,[8���ed�oC_�e�f9r����iޟ{C�������%^M=u�4F�x���,DG����qK*��L��C'~OA6q1z��ކD�n�g�r*4����f6�Z�Wʔ. 4�s��^:��{����H�����2	E�����2�����nuuR^��H�O�3
h��3-�^�l�ȏL�D@��whYZ���Ip5�u�KT��3yTљ�^)o���i�Y7k�+��k�*������?��M�bԛ"+:혞[y ���*��WNHgX��
}���8�p�����Z�R���U�W��#O�A`��:��T�GM��W�|$��qN�N���y�y����g�=�֧��JsH`|L�,�Ty��a]֞Ĵ��~�M�\���>S�,���)����)������Z�̂=��b�
	�|'�q_ԾE���~���m��\)*^��Xu;֊ʳ�v6$�Z��|�¡3l�ړo�m�["eg~��'{����;�1��a�0�?Xh�Ռ�Y����`Z�!�K#�z�u�ju����ѐ�@#G�-.�j2�(����N.Nv����yp9_���TcH��ùߞj�t�t(�v0f��/��+�@��8&Cc	&�!��+�!��m���ƌ��3�ok/pW���"�d�[�0�l�m�d��iCbRz�I�ٸ�3��ZCr���N����
�L�h�k��b��T��z�m*y��Fʹ:)���m./Qq��钊mƏ��&�%��I�ڦKB�ɏ�kZ���5t)udL�t��l�n�O䊴�u�7L������x�U�l�gc�����>�)hNUn��Hq`�d��Ża�,��+�y�N�Da���y�n�/%���z�n6?m������!�ͨ|X���䃱�7v恇M�c�Q�k@�O���;EѷJ�OJ���&��C����7����%Jm�w\�9�g�,m��n�ލ�U�������>��8{�Okk	����TP���joP(ŉ��m�f��7\�z�� �+��ϫ��"L��Mnj&���	Ҙ�E��J'���Ub�5���0�ԑձ;rvm\F����/�׿���o\T%-��?�(�3�g⌫����P��
Pj��oY;��ˮ�S����ƴ�,����;6�Pmz�)��Ƽ�6��v'(H�y���2'=���jZ��Z��PoI ɆԌ�1�KQ}�S	�Y�������j�&�$��%��M����j �cܑE3un��~�]6_6��n�@�9i����OȤ&����)�?�w���޸I&�)>��l͗�]�:��UYp��cв��6l�)�3�$�~ժ0Xr�m�n]$�����!�D����I�/�@v7���V��wR��/��������~�`���K�g�y	�Ψ�8��a��S��x����:�+P�����#KDм"�_��Z������a��?�!�?E���.$[ɦo��0G�s��ͅ��l(�B�CB*![z����/��`2V�����p�E!	�@��8vE�$ ��igjn��Ϡ��Or�)���dX�B�v�x5r�n��R9�T��������C��=c�������W	��3�')�=0,���3�hౡ�6�s�u�D��(��[6�%+��"�q��d�ѵ�N��P+���
��v:'�� �(9NJ�¨ކv�9SU5��F0��K��-�c�V���-��BmjI�s�ekϒ��|�����3xu��[.���S��k(���bS���l:��aXC������A�}�r�L$�>:�E{5[���Z���40���?K�� �.���U��=�%#J�"2�ϩ����Uo��\fm�`�"V͉]����]� oM����P��W������d��gɀ��Z����"�1.����Zr[;���i�}#�!���{u6A$9�٤*�j{�Ã���:��!�ۉ៼f�55��Iۡ�w�ݱ�{ƽ��O�Nƽ�!�,�.fO�ܶt(Xzm�M�'<��ES;�gg��*�O҆.?�7{ ��&���	��mW�jD�-��Ixټt�:�HA��ّ��{V!��:
�	7�d�zc�u�'�>�����ǰ��j�"�~���~��^��S5wW�cȚc�$
�<�u�驐��qn�y�Q��<~ś߄�1d�L�aP����aF�Jq:��jL�u�-��t�r��eJf�`dͦO���:���R��0X�N�*����i�8
�!Do�)�~?Ѝ��9F�)��l��t�b�p�z=V]~�V�#4���W�&��p"�*�S�(���a�WS!;nP�GX~hEm��b�/`��8��4�����-I1oG��=�z����^�_6 �j��vt���f��+�X�\��CRj�jtd1�X���������Da�mطmY�4��j��~���Hi�z�Y��1a
$��QHn���E��m�&P�̕ ^u;�r~�`AO�|���q�H��0����!�
��i3�4�>b\qingt_�`-��)�ӛh�/��:������\�Ϙ��Q�1$]�mt�E�����uf"p%s``���~�l���!�H��muV�9��u����]$���m|.`7ϻ:��ͯ�KC+]h��	O'"�}nϒ�U�ϡzH/��[�tX>\��V�~W�:Z�
�Ȧy?|��'2��]6 %��.��eu{8��5y�dE�\&��!�����U�[S�!WK��y��@x�<�EK�c��}8�������{4�W���MP8��L��&��U�X�O�|K )�x�e��J�r�_tB����Ƙ�$-����;�l�N�L�K
2���7�O䉥Hrcd��\�4.9�:���Ni<H|ԃxg�\2����*�C~:R�5�:��
�yԮy�mN�,��5A��e��P�SM_���=�E��@��D����w����Q�w��<�|�#v2�<���c�)�O���g�>���0/�/cw �52��h`[f�����T�}�ip�"��<����C��r�x�H��NrK#;���w�����e���>�4P�fFu�e�@q�\�z�S�.�_�>2?�w!��G�4�h��_n�Y��>0��r��P8�`��$��R/��h�g�/�M+LB�!���7$ ��-�&?	�<y/oh�HJ`Ӧʎ�|��h�.Z�7w��Α��]�Q`a���	�+V�C���o��������S(c�
j���@RP{K2i=\L��hk�Ԍ�~��q
���m����wQ�!�Z�.����L�D߽&����y��C|V���͈�Հ?5<��$�@-��ù����) �]�@%�A��\�Q���r�Lb�͊�s�Z���^��a��~�K��J]��-vl��TڗV�.4������ln6ѵs�&����:n���, ���[��<B�K<�	��fqǢ�i(o��6� C�A�����Wk8�Vcn���v��"��[�>�!rF5���5Jp���[�M�!���i��ve�UX8-�u}�'y��7n�[Zd
S�KM�'�7�i0W��-D�5�ɣH���Hpז ���x�m;[X[�*�Ps��杮����)>�_��X¡Ռ��Ο4���?��#�=E���[u{�����)��#U;[���=�
�������sY(Z<i��8h �l�- �I���[�6��ƕ<� &R`��S/��>P�1F��_)ڪ5J:�~�]x!�Y�bə/���q�ƱQ���#h�2Z+k��}����
��X��s���Z��[:�p]�x�O�J�4O�	0��Ɂ�����㣚��GU;(�4	w���A�ɨ˂;�Iȼ'p�5e��޿�T*����?��S; ��y�7�[�Ø,͑�JW܅��Y�U�&�lL�b�v�.6��+�܎�?2��Bǃ�}���Zk�)$�mh���eQ���_�E�r��S�n]"�{pW:
m�6��$���+��;c*�>�Q�L���n>�`5��%(��Bk�Ų�:�[j%`;�g��1%/tl��W�y=��y�.���91$��&�;ޘ5p��v�A���F���`�#��Dٯ�$���`�e�zH&�_еq���`,A�fY�U
�����.@�̅�Ud����7c�(��������5���j�~pK>)E&jt#	éoz��ґ&:\��;��O�(�u7�J/�]�=�(5-���l&��(b|��a*>��_��L�qE8u2�%N�*#S���ƤC3��H�5�]%7��	�|�*hQ G�oed$s���n[>��`S*Z`��U�*÷�_h���1�+#ɻqF�|�ƕ��㋰�����;��Q�|kI�͚ŋ�+���;s��j>]��S\��TD=���fQ�����S�O���&[N�']M�&�
V�&��i+��i�	*��5ڑ&��GYW�§Ń�M
)I��1G'�� ��l��;�7�����k�>h��@�V������G$ wS��7�Ɖ����ʻJ����ǹDf�yzԽ&U�#?��y'������LMtz:b�R�.w�s��z'`ZЦ���|�q�z� 0e˖��,1�^|��4�G�F���y@��g|�9�0�3ޞ���d�U�"�Z)X��I�)�::�tP6�aH������7���EN�o��	���$hDPm�	��fP���Z8l|�i��_��N�>Xr�i	$o��4���W#�k�����N��*�����c�����L�SP���m�s�%M��_ƛ�}7���{,oI~S�#QWt��(����%���������y ��*`&t�2�3�e�6g��Å`�YTS��������=ՅDP׿��lh��?��aT8)]�.2��D���g��m�����Q��VG5��9d v�P�ZLk��je����g7�R�(X�P�2v~�����J��)�U���6F,>������/�NӚ;OԽ79g����٥m�΀����^ϒ�I��Q��� �5Q�:T�?$�����m����O�F>�P�,� ����5�!�Y�)LxN<d�r�r���Z-��pP��4q��Jv��^w��Ƚ2Ce����ᜉ�
��Uu�:5��ۋ�|��f(}�����xbQ��Ҧ.ې�������E1c`��� ]QV"�C)s�ܲ(�y���-]� �¤7�.��g��i
}�{�#C�[TT�\D�`lmP�ү^�N�ga�a!�9�-ne'Ka��j����"����`�[����0�#oA\_v�n�Pc6����Ʃ��G>����ݬ-jNƹE���S �B��<��w+5-[vq=V[�O}�B�No�{ʕ`����Q����Q0�T�k�)2�EW[T��5]�t���a�"��1ۧ�_|�5S��0�X&��$י	���B}m�� �� �j�I��~Kw����BV4��l���fQ�v���.���H�����j�
�f��a^��ϵ0R"pk��&�����?�.���Dv3�A����>p�y��8�z:\��P��=a�����@t�앦�[KdJc�v�Q��BA��_���bF΀�҆0�5\���5@��[F L8m�i��R}|������9�n|vOMR� ��0�޵i�"F�4����A�J��G�J�Db��x��N��r�o6<����Em&��ԧ�Ztϙ4aDB��gW@B� L�_���쒶=�0`1�FF/?�zG���><ͳ���6�^��P}֞3�R"�٬V�q�V�{��/L���HŷI4�� ��R�΃XYT?p')P�E��#���8����{(s��`�%���qhY<�-��O,�{���d�����ud50|@�ϴ�~���Zx�����r�6	�ԕD���O��ǉ
��?d��� s�4f,tN��V�lqX���=�&�E�B�Z�:�#U���U_�#u��04i<̨�T���͕4!�x(���b5���zK�_9�m�P�i�.�����c��=����J����:�Qܩ��%K�?��]&l��YTf��k�.
I�����i��9�z����l��򝖤��c���n�8�C<����6�4�qhO�%^�4yZ<cJ�E	Y���>wqa��a�=�i��m~���'���0B/�u�$ Q�$������I�]v �)��#� L8K�;�c�s�F��������<�y�{�G%P���cͳy��]� <���*M<a彆ީ��	s�������=�8��N��R4*�֟��)ʏhlW��*�*��Onj��!4VJB�P]Dt��';��^;
�\��]��$��UsG��q3��f�Ä���:=�������[u���J5칬��Vӵ:�C(+��<�^������77���Չ��a�޶ͣjB�p�Y�p�g%���l+�+g ����m<.��0S��n�
�x��H�-����J���\CP+����UD�����<��ڪ�w��X��W�~'��T;C�CtS�/V*V<��S)���re�ނ��09ݢ��ƕl�V�ln��{�y� 9�
�Ԯ1�TP4 Eq�|͘�g���D����h���w�+'�3`�/±A��Ƕ#�&'##�]0�����Wx�;SU_"���,LԚ��m�%��b� �6'�p����!͢"�S[�-�" ,���h�f��w���#���9I�ӆd�;�&��X���Q@����I�)mY8��r/�l0�>��g�i���ʲ��u.�P� ��e��p�����>Kt
K�*�u�\{v�y�'���K TCn@AIC�#]��i7<��l#>+s� �>���t4�ǅٞl֌G�U��w=jWg޻�X �|$���0����98X��R�'18{(͞2ie�Ӵ}�O�G��XAJ������q�T��m�͊�ջ�����ν�e�$�y��g���n����~=�1��5ޟ�삑�NĚ�5J1ʹ⼴�k�Uk��r�&7O��x;O�� x��j�Z�J.����d��K��ʂ/F����،�����b}���=�2�p�N��K�bȃ��8-8]J��w��!L�2�[M'Or��W���H�W2 6~�$���"�w]7*��\+�>@[r�}�PX���tp������Ev�Y�;Y�E���r��+�]� ���'v�ﾯq���6v$������;	{s�0u1�
=&�d�1'�I!OՄ�Z��_^�'[W�K�?R&
�a��Tk�>3�1&�/�5��R8W�>�:�8�}A���ZuH� ���t���)K��oF�,59�Tme�9����+FWH[>|��~�o�-pBu����c]@�Гj���b�!����1�X�R���	`͖+�p����E����4uuT�Q��Է�_���!��p�� aR:����s����V�o��A'��6��ϷSn���>`9_��D�Y"����ת��s�Cۣ�1��8�0B��گ���,	�1�K�9)���qi6$fk$c�j���!���0��JY*z�*@.�f'�,i�̘�A�=��|�̓���H������V� TԵQǖ
�����xf}������'[��T�EE+���>a��[��s��8H࢜����)bP�,�LC
d�W�R,����Z�
揙S�8�%&tS4t�QG������6{?���9�%8ޖ{�N�*��(��S���	vc�xFX�p�+|�,lଶb�o��8[GG ��\����y0�^��/?H� !�
�ώ�˂����@;2C%_�T6	��޸�n��]Ռ���;?z^%/o����߆�}�=����k�>+�WW��l�5��!�s���$�(TU!"�����I;-���ʎ'RI����%��6pb&�S��fU�&��ï��"/�EQ�U�ٝ�
���>!�����7�q�/ i�"Ͳ-�&m@�*���^+���)��]�@t��~�wd�����γ�I��H�>]j��I�/�X���f
�,$m��`H�Bp��˨�Ys�^qش����{^$8P�	��aS�k��p[�K�������ׂM֨��z�2l���'�_3�=�N
j�o�[��D���XĮ�(��f�j��b3ܑ�������͔2]���E]X�&�5<�s�b� ��� ��AKtn��T3���No��Eb����4xD���Y�|�T��fZv�`-��u�\��	�ӿ���i�j�~��i��1Q+Jy/��gi�n�x9ɹw#i[�0����-q���t[�e��ּ��"=��ŗa
�I�Z!�h�J�e Mm�҄��1x�����*�A�����8S
-�����d=����XwDˌCo���Q�߉��&}�ݫ���Y�Q�-���G��AJj�K���M��'�{��⼇��������v��O$��5)(S�V�ú��F#����8%u�Mi�Kdd#70�U�=��� jg3�����r����Xa���ѷ�ݔO�1V���+�g^�C( �����r���k��|���M����w��Qe��@/��� ����z�h����:u�֮����eH�P�@t��qH�:Y��Ƭ"���xD$�YA�J�
���8��C�JԖcX=��.P��b��#%���p�|�>�	�I�h,6Z�ng����h|�A�-2��_����E�*��Z&�?@�j2�T��u���̀>��DEeeC���w��c|l�5f5��pM��E�p�o�F�;\Ub��os�|K)���o��(�I"kc\�H�����2�6C�;V,kl��b�����������(��hISE���Aƞ�b�s�
���#�YV�-:LQ��n������-�����J9������*���( 4�w�UZ	!�s2p��N{�;���B�Cėu�R���a�$�9�#���t�G��V� �n��v5�����	]�d��q�P�ﳤ~��*�}q�����%[��"��fzO~$K��E�MH�b/�sO���h�}M�H�I���<&1�PX��-�I�עF���	�Z]U�[pq)���?����g쌒������۔um��%���;hC�;�f=����kC�<c�=�CV�t+�v>$���h;sI�~ �('O��Cs��ٗP}�$���j��nM5<o0�.�j8;2��X�I��X�CK�t2����_2�)Ƨ�"�7������iv��07Z%f���%ۓ
i��ob��=}��T:P�ǵx�&�K��}��)��6��!L�H�Ir�H����]!S��\So0�n�5Z�R�qF�&�~���p�yb��Y����K�.p�C�.F��vنJ�f�`����-/�'K��f`���U(��
�<w�A��2u��)>.:혬�(������v\����[��5�V["��3������(�uIc�T�7��T�Π>�x�8���%k�f	����"]��׳m������ߓ�����o��U���a���	�����y?,{v�y�����s�8�Y�A�7�Pz���vF�{b~3��A�HLGJ�-��|�gl��)�l2U���Tl�7��������tz�S`1NԀI+g�xt�ʬrv!ڊ�����#��
);".��("�E�h
��5X}�=O@y���J��z��N�����,i&��	 �'+ɉ^�տ�t ���J�ѫԁ�~y�K[�&l�C�3��T'�\O�i��ɝ���2�69��D�=wJAt���4Y}�I'C��1��%΀��t3l<��Ї�
	�3�*���
9�E���XH5z6c��&]hsuf~�Z��a��Q�ʞR<�:x1J���*����� X���9rU�9y��R<�<P�'<B�М ��O�Y��i"��˩��Jn�&!��L�ɦ*jҕʾS!ppI����o7Hd�J��F�oS?��9@y\,�_��B:��oUlwW���Rʝ����U�fѴ�$2��w�nׇ�&�.�)��J�@GI�u'w�f$D��E�^�1K����Tz�_�@}ɉ�_��m��袅Q��7�6�O�1KIMs�ނLS��/g4gx���zY�p~.����8���Ԗ!�q.��X!�R�Y��]\ �(����=/�C��d -8:����˹;}��r���_�[襥�
��F�l�?�����:�������o��!h!���a�pK,Y��g�84+���{�)�y'7ʬ.�_X�F�ǧ�Uh:Y�?����{�����h��&e���"b��P�U���NW�����>{ᐩ]��9+l�yR��Ot���!n��UM�T�t�(]Q���|�'@�l�Kv�0YU	<��Z�̺�K���q5��W=v�=��-ӆ�}ʆ��J�D9)1�Y���V��f�]D��h=��|��P����R���@Ȓo>�N=hl��H�Gb�T\�����~ڊ�c�sELc�>tq->f�����A�����̍�_��]������!��j
�pF/$�C�jfmڢ�Ȍq��-�I��8r>PȦ,�I W�
h�����c�s?B��>p1�����o���:X����󦲁�����%q����oz���Ӗ�ʐ�g���|9m|��L�^ 	�'9��o3����x��v���^Ae8��}�J
�<ɮ#űp*���9��:�$0{!�5�N�=p�=�����n(=9b�Q�b��l���I�H�w���5,�-�ʾ��j���^{N`?���q��m�	��6��~�M��X[�_�E��[AP4�{�����,���=�$༷1�̶]��3�ނ�?��x;��d�$�2�Z����[�svDՙzHz����:{r9L"w���RWn��[�ǬȻtf��S�D*�ޕ�F�b	�ܪ^zi:��NɝM��Y'�{&��P�ҵk�d1y�.�ԫ�BOxC���m�Uw��
أo��;,7P�@�����R��;��7߻\���Z�Q���ґ��)qp�?�tm��D�w��:���=�)m,���"ଵ&��J%S��7�z�Y��U e6���c�)�~8�隌��&����ⱖN7�:����ר0�UPG�ڄt�U��H���U�ק�e|<t��;)�f2�iVu/Pzu+���H\�ih�)�~ ���<
[��ſ���yq�|�?�1l�,X�����OhPs��Nh�*I|"[ౣ>�$e��m$1�<7����.�'��ߑlL8&%�J^	��3�����͐ E�� B�1���i���m)ʯ3������T��?n��[E�>&����#�6�}3o(#��Mg�%�F�C���&>�9�!>�~����id%DI��^���<x�"���┓��d���{k���s��P��l�/�����h#�}�C�,�)��o����i��TP4T����|�t̙�p�v�X,�k�Y�3�:~�8��h��<�T�#Q�,\�|I���EP��?_�$�tCN�.�����C2��� P�m�ǭ��VTȓ��I�YQg����I��y�Z�Yg��:[�l�FI�r�o�KC:՟lhLgnۤϤ!������T��Y����B��8p	���T*�!��EH� ������C00F)��-�$��;��IpX�=�����c�}��p��ic�<}@��}Z��n��\�D�`�T�:���}P���tH9�3� eJ�p	"�:�@z����mN.�h[x&��-��|� �_��@�+oʳ��Bp����-�9XIVGW�K�\����5�S�^fW���[��W����&�T�z�(0�/0��5c���o	(>C���?PKw�uu�]4`��T��^��M��G�sR��Ӈ'H�7�[f�[:��)�����I�mb�� 5�i�~�5�tK����Y�[�i��������	�̺����Ͼ>�{6� r�-�wa(����[��jAD N(���zA=�^�඼�� y����ny)0�Y�?��o0�S��w�O����z��~T�"�L-4���q���I�~�(s�����,��8�1M|���Z�j��ȴFz�>�D7�"|�:[b}��S7��W�mlmq����9�y��$մ�&��bN �ȷ�z?4��z�0G_ۻ{�]����
�:�5��������&i���!�I����)Y�\�6]�=-�`����Jmݺ��L��Yش�5K�����*� D���N�m���F�!�l�I� ��`L��0�;V��e.;t����� ��/<C�#�`�	��Z�&��Hn�i�<���V��{�t�q��v�#t�n\�Q��Ä����%��\0�F���;�1G�����!��Ǣ`�����Tk�Z "vTiu�0�hB��#6)�Q��p�r�_���+�����c��\�\����ڿu������L�8�2c��ǻ~,z[���\�z��M��bfↈ�(�"��O�����,��f|��ǣ��i>|"�����*��
����S���!�[oL�}'!O��U�*�ip��k�<����6��g�bc�u�s�6�?��.�k������K>�0�� W~�N���tC�&����0|��L���rX|�n%�f��[I�4H<N;@rq��q��>�S��?1I* W��~��(@R2���Ws~Rr۸�Zѻ���@E�;RwtW+=󬀳����QE�ΰOa��i��q�Ѧ�K4X���#���|��B��7�x�T��)�H@����Q���3��d�]}��F<��'�Le\��!c��	��6�SH� �§��g��O2�$�ů��t����&���n���Wf��� �rc�
-ޔq�>nE4wt���wkk(
�jp拫�"��Ŕ��bD�Y�gӺ�VƜ�h������4�5��sN��F�^���C^��3�&��pp!���uBR+p|^/e��/�"�>��3���Sڻ(S'ZZ�8İ�>$�����k8������e������L����b��b���7�a�#Z�DG�u������$�^��C4},��̓S�3�\0�A*3?]�ٰ���[��W�ep�v�Ҧ
�2x��uv�Y��y�{��l`cM����zةe�Wl��$::�)`�lpX�D��R�@fj�SDQUStܖ��Qt�M��u匏ǵ����p�z�A��ڊ� E���E����ǻ��݊
�m6�q�E��բ$n%��ZM�~&ycXDW?R8E�7i�J���{9�0!!U�X��B�Ӈ!�������2��������<[I_Hq�{ŀ	^t��9
��;4q�)�J��"� ��f�.Z>4��R$��zűk��V��/���87�n9��Pɹf��{�`�\����7Q��h<���iGE�E?5r�X��FY���[���X�� {�\���h��еHP"@��*G�I��T�l�$�w����+]5M��h���C���\�ٖ�<^�ه�(�;�����������^{O�un!�t�.�(�)��j��D�/tJG!��ͷ`�~�4�8 >�&������d^�A�L��^�t�d�ij�UC/q\|!J�7��!�"�wڒ��S��,n���O�I���):L�����
D�l"�p�r��-�̐N-ߠǄG
�E��4j���#��>u���gڋTo������O���u��V�o"Ǌ�R�Q��q\��v�ߩ�e��8���b�Qͦ���ב��|�����=6�~岐�4��y�4��b��X���K��8�H2�D�$�<8����t+�v1��?􀻟������ٻj�#X(�-�t�+�b{�1�ݦ�=�g̳O�r���y��{��]lZSXC�;!B��pno��=i�o�RZ)`���,X,���[�LHq �A)����CQ��p� �Cu��/?�����eF�i�/�ْ�m8�{a���f�&�v�K&�T{8��j<�$x��ww���S��鮏o��M���y�so�tB����_�-<W6m���A�����s꟪x�v#Y�*�����ٕs���`?�9�� ����2r���
�e���5�֒�5F�agE���Y����E5f��ӵ `�+q��:�F�K���X�'��B��~K�����P	|7�+f��}�q�u��:-�Y�ߖ/�
� �?��7Wx�p/F���f�vM#���:WI
j�ʪH\�:�Y�%+a�w����4�����ʵ|��� ��> &���,g�m�19ʎW�w�a�xA�S�m\oO���|ǁF��`��F��Ig����B��:��k� �䫑j�Yx��C�����rK�� �o=َf_<c�u��R�8�n� �c(�)�@�?뷪�L]�ѳ���r'ɹ����`IM�'�]�� ud��8�}38���ܑD���}1DOy'5�d�����V:�g������	S+�����>ac�I�"�<�M����V��:QkP��$�)7������G�!q?��
dFu&�i���^8�H�u_{�s9x	G���8�F��y�<(n9����<C� ��
3fŷewPe��{'X��>���)�V�"N<�Lum
�3o��d2G��4:"[6�4D#���Iџ�ߞ)��a�"z��5X��1L� ��q&Q]\�&7�У	:2�'�\�����g3���9��d��P4WKĉZ� �=G�朒F�р����v��}R
��iש�g|��~�`lK������o.Z�WW������+�Q�]t��jV�������:Fl�Y����#.�!���Qp��Wtܨ�܍��AI�4�a���#t��0Zg!4y9�:��=>]1!_^��P&_�`�Z',��L�o�B9��g��-؍~_��Q���>�	�Y������B���8�X����â��y�,��31��q��D��BUc��C$�U�RqI�0.��m�&,h9G&���3 1��v����?���~�}���8�;�H�r��D�ê�´�����YKE~c�0���#�ه�O �d�d�g��}g<H����xǮ�1e$����-*S����U������!D���bW�8�+��F� ��'$*S߂9�f��B|�җE��4�"8���qcӤC�����g+��Y}�4cjg�	��;���V��S�|���uq����v%J�94e6/�_vVA���N�נ�;j2�|��m3���$��ͱ��^,��
q��*NHJ�O� od-zsr��f�$��>vk"D�)����5H�h�Ћ�O�~��#k�i��C2�}ik¸v�p�	�c�<B	�`���9�����9ɨT�'�;L_���&��F�qX�������iM8�h�g�J2YU��I����������.�u��ُU`�e��-0��[��d9S��fځT��2��	��`��F�S&��f��9�X�Y��|W+`T�@��>�s'jM;jC�Hq=M``,��?9۲�nٌ�n綏����W��0��*-���$R�t��,3��&��A䟺�O	���*d�m�*1�Ӄ��@/�X�%�]JC�x���_�Y,�cz��0���!_� �ƌ�$�� �T�K��l`H�&Z�]���@0xG����Ux`���s.����ueEA���%<���C8����'�檟� ����A���F�{#?�$_���5�4�v`��2��2]��2D.KZ��38���$�õ�dc���3���m%��t�Qkʠٱ{��B�I��5C�9���*,Mib
��������a�����lh ~�ԕN�Y� A�?r�%�/.�_N6+�p7�|�g�ǥړ;6��;�?�?���[��k�Nս���I�ML
��EU����g��0�*߳�Ei�W9e4%@HԹ\�ڷu!c������T��4��9��u9��}��������.z�^n8 �^*�;,�EF��&�=�>�n�HT���0��`h�a�f����J�~���;�$��nT˾�p��U-���	͸Ï�j7h���)�ql����"��v�xEԧ��n[�]R���,uu���V���'��9���x`��]�s�ds��ޑ���!0�T�+݅D���Ӊ�|���z48��!q�������Px1*�� 6��+A-�^%Ә�*
�bۇ��Æ��5��aAS�q���}�Vq<K:p�K2�vˈ���"Z�;�՝��@uJ�<�ѩ�j��ʊ���T��[<S�8L��f�Y=i��]<Oێц�
��S��OJ<ē�m�6��31��z�U9�R��_m=4���V.*i�}�K�g��N,cnb?;|^�:�����7T�U%�k�v���M�?[{K��qr6�wƎ���������1#��F2*5����P�n��^�Gc�j]���'�,�|��*J��A�!wrЯ��!IX<�s��F`G� �)�F���>H6�9R�Be,���cu+��4�s�:�\GVx�~M��>q��Mp�����\Vt��2�ֹ��A�� �OԡGź��Y�t_Ht�s��F��dh�p�X ��Hs4�v�Za�fҥ�ے
�ޘ�-[=�"�R���(>�VXW?$ ����LP��[��(�U�`��OOs^o?��UM�VN)� �l�-qO �n��r-wڵ��#�� �U� �fmN<EY��A/˄Y������=����s���ؽ�[5
 ���E� �����+���9ZmiT[M�9��D�_m�ƃ�E��E�3b{�$���)t�L]�Y�V!~�-�U�B��"���0����V)��b5�*��֪��@pm��o}#)���r9��ळ�D�	�k�8_���YG���mR^F�T���fČS�g�~���G7Z��i�@��*�=�^�yYt��`X��P�_�	!uw�"�`�[�l2H�>*��=�l*��Lw�}��#�6h��G����O��5R��b� t��� ���Jk*; |F�Q`t)�)d���9ҳ�?L(qM�A��+�q��;\� �7k�F'I�T�dY+FP\����ؔ3�}~,M�FF<����ӣo�j5@c�*��6j�ZT�4U׬�h�!��{�AfS.�/}=�b����|8;�C��m��j�dc����zu�3E�X�*��w*Iَ�#[c':|���	**�f��IO<�?�������2�΅�a_�N�
�l�N����lO�6�ɯxx��і:���(K*�g�z]���Q�.�n����p2��I .Q��5p$s������	�ePۚ-ʻQ�=	E�Dy��öVHԭ;�"Fu�_]؎�Z�ED$Yčѓ{~��o�W��~�Ǹe?�ʑ 2'ԭ"X�6E�;ås�̯|�ؕ&"�`� � x��8�Ԙq�ܮ(�QB�{�-8��
��aOGub��l?N�cH�)�o���O*6hjn�$�n�`-����qȊ��$��;G�:t�#��df�@��`�p����+��L��C˸C���GOG*�#Ŭ�%B�)k /8X�N+;�z����� QM�����J�6��®��*|	a�6�T.�r�нǴ;,ץ�8ɍܟ���8�ny���|:�k��?E�$7P����o���J]�ѯm���ځ~�yɆW�qM�d*�Q3��P���z�叠na}��:���%0JuXy��5��`���ts踮M��vv�5M�4�T?��32�EG�l��b$���a�����[uN���M�ը�d��#E�-e�m]�DMs(!@z��Z���b�����.�`�NY�w������T�/�1�)-\)��I����-i?Ur\�-r{��6� g5؜冻��Hg�g�_���E����I4�Jq:�
pN�x$������b��(�#0K:%�}�~�ә�>,���a��[Y��smw3a9Ҷ�_�)$M��Mx���ٽ�\��cMB�.Th��@ �����R�`�p�u(r/��s7*�SQгľ91��n�fR˹�5�XE%�Y�o������Ds\FXw͈�q^υ-Y+N�Z�1�eɼQgp���E�Ҕb�`F��k�Vg�݆��t?��A�|.�]P�g����@�xRB�wSqZhvF�����0��<��;+��l�@Z_��>X����q���(8��4w��
�J%a�x$γ�@X��5�v�Vc�e�y�$�=��(?
�g����T�zQ���\L�A���Q?1
�ɰ�T&n�X<�#�S�>4*��7ᨯ��y�l{ko��T�V�l�Q��r�EK��V���FJZ]�8mhB���D�*��U�9Ե,^�	2�P�_-�pAl����m������ⲽ�[�w��nL��#Ż�����p�K	��)�nKD�z�YR�^%(� ���1�Ғn�}c	-Q�V����D�l#��}%�6J�� m�ͽ�]�����r�M^��T�!���phϹz�F=9D�rh{B�)��w�v��k�\��ߥ��!���������P�檠pA-jt���$+�v���_��3��-+K�=g��x3_��U:�C�u&;�7����f��
� �%�_�z����]�\��cҊa�,�2?r*�s�6�@G��do^��9#�h��9���p4Y�ڊ�a\�� ��9BE�UɎ���gwG�#�L�zb���2s��F��ɵ�t�.%.~����l%A�X(�p�ݚ�N��3b�8c��a��b�|p#��G)-����,�y!4d��6�K�+�ō+��@C�y�e'd���|����|z+*$���x���t��\z��`3��i�~9����,�K�]��Ø�c�ZD����Do_ �#_V��s�y��V]�h��_Ϣ�\1�lY�(��O�P��}T�{���E�F:�£.D�����T�fn9��ԕ-5�[�d�:KL�g3�`򆚁�BJ��WV� �N��;0��h���"л�z�~4�P�����_�J;'�[Y�/��[Bt=�����7w�oIL�M����s���1{� [S�k�^މ�^C�����aW`��5�L�֝- j��;,f���LJ)E�Z�p��[��)/���u��m�8���m9�T�Hf <Q�R����O��Z�VG4̭yG����`�t:�P����]���\Ɩ�^�JmqP��)�jCw�����$��VƷ�q����7*�$v�o1�1џO��鉔��Ӷ�j�JI����jI�yq*H:�0�eo5&�$�j&�PO ���*(���������T���g�̍�⦢e�<�d�>��V��H5]闤}e����?��)ʑ�SZM��r��#>��) O��l��dײk|W7.���Ù�j��OV#J̌٧�RV$]`��Z;K���K�4��ā(^��+�����7 f�*���[a��P�1�^۔��TDئ{Wm�1#�#̹�цJ���'��E���p�b�O8IKI�n�������l���������?�u6&k.�k�\��yaɲ���ۅ����%k��^���$>�B�G��w�-�b��PM�{�X�uZ'Y��Ta'�v��]/�p[ɝ擝R����fT*T#�<���$/��%��(kV'�E��s��e���������h�Xo~T��I�=�iW�=n:�������4(e���PHMȷ<,õ����'�NS1�ez3�f'j��E����ʘeI6�����m%�qXQ���|�e0k��6��6��M*���RI�Bd,k�5��?w���KTjk>i%cKO �83��@��cSc�p� ��YX�������crdQ�tS��լ`-lQ�e��B��LV���}sܧ(�*���k���<26 �#�q�de*�W�F|��#��T.j�u�R�ꓶ�~��L1?�*���Z:���B��n��_�<#��y��B4�����ɇ�t��r��e���_��d��9�����~;l�UH�g���:�O���,N��y�EHO�j@����K�O��GV.�tQN/e���؃Aۆ�Q$׏ȫg��A�l���6�DI��Y�\9n�*.r*�k���u�܄&#�@��UI���M��=i�?���L/�3Ck]g8i3��N���X:{��"`��^H����R�F޶S�6D}v���c;�X;t&��gi��Bz�B����Q�ql/]�k����I��K�?f�f5d��z��y��WM���]��j���SW%�5E=&`����STz���eep�f��:YLay3���`l"���4�q9�����1�4Ƹ��P⍲���qr!�kL�$�Iy������ ��}6�O$(�5$
.��gG�U�����wֶ��GɎ�8�99A���37��#�w`��E��u��Ԙ�_|��'���H�W��Fyf�[���_yċ��g���u��gx6xm��xl�4�_� �T �h�׫��["�I�f���a��N�(���6������ӺU�1�ؙ��}�h�0J ;v>�Ȫ�S���U���V�秳��a�dv����U`�t�.h%H��8LW�,m=�c~f��߈p����1a�S�ú����K�iKs�9�]�`8�X��0��5����'�z�-�C�]�
�����b�<����-R���g]�۝2�1 �9жU������9׫����G�	L�x�~��Q�CG���6U�q_��:����ŻGw�-������BG`M�A��Qgo������鐨J��^��B�6�v��
yd���CC3��Ҟ�ʏw�(��n*Ko;ipIaTl�>�.�ʀÍZb�r�ۭ���w)(pXb�i��T�i���9Md)��� ~�P�;�$5�w�KH�ے���z��ׯ0���ա�#;\�q3ٚ�(]�O���q^=f���a�t���FQ������G6k�#�RM��x*v���o��-���?�%��	��y_���<,�lS�fΫu³dh�������11��"���2oէ���_�}��~R�f���]�&/{S�����4W��V�Ꜻ"��A����DJi�%����1F)�I�����oz��@i�R�%�\��`��3�X�Bݵ5A8mM��v3j�v�&:�~ՠ2'�� ��
)Z�Ql���3k��ɧTs�~p�n�zs�,o��&���7���i�j�>��-j���3�o5����� 2}�=���0��������r�|K��#��(C�)Qasr.R~F�,�^C3��_�kWsa.��~x�@[L%��c��߻&�l����^>5���fg�^��װ�AP�M�بmw�Z�b:>��ӽ�	���N�~�ш�
��?L���oX$M6����4�)�W?��H��ß�<��O㔏ū��8�)J&�������w�k�?o��{�m G�[��~,�*����8��|!G��6��!vj�",z�>5cRk��޺��������4�������K�en�k������߂�ٹ�6U��"�x�$�_��Ү�I��(	��^؈��{�B&���vE�cƀȗ��Ѵ�1M#pF���v�݇�Uƌ_m`;�b��[h*:�Z[K+�����JZ�1:Q�JR�����I<�������D55��;��&|q3��򼴄Fz�'�t�����"�6����L��"�� ���t*m�����q��;�sd�D��S�ә�0���T�(S�hJV���˚�����ex�2��ֳ�v��eT��38֏0)����6�}1ב�:Zʎ�AS�;�s�
}�!��N|�[��u���֟�:w�ؕi5�f&�S}��&?g�-1�B���Zu�\U�S����܃�r�mr�t��Rm�s8gj��g�p�(C�ж#�iHFp��,fLr�]G�)
���̨���qo���,��h�[�%�Nn�5�hX� /;�:
�Nr�IgU(U��8���ft\�h>�&�Z�a�?Ex닔#��]������"�Cwt���MS~�tV�GF������O-RQ)!�z�$
�V�;R��ȋ��e�����1�Q�hJ~9܎M#����r��Q�h��`�C��ij��ܘʜO/��%mאw�3u����Wz��>H�`�	}�zT�+�<�~	��� ���qB,��c��/��ߊ��O)���0���FӤP�1�tΙ���6���Ŵ��e�qG�jwE��֦ܮNGb����De��4�A"U�g����ܹ-]�C�y�&�����y�y��2�\��˻@���jR��KFR :��u������	�� 1\�׊���)+���3v�
K%�Q| V^�n�5��xֈ�!e h�w�I|�b��G6��o�׶�ND���B�kR��z��ѻ��P����X��@�_�f�9� W���Q5+*$֍g_��:텮>Ǎm]m��I��`�/T?���a%K�~<<� 7�F�d?z�^Mޯ��+[a�$�Ӌ�
^���駹�YS��R��� ��Hpr�Ge���(��A)�>֊���Yzn�� �k\��/-�s�����{��>c�п�];m싗`�*����b@+b�I�
��Klx�X@�P��4Qp�.�dm�.�J����u��N<�Zk����nV/�q� �w��^��WKK �y��af9a=v�G��[�\�Y�Y�O�/�|ۉ�2n܌ڒO�jE	��q�	>E���I6��v�,������ꑎ+����ᕳ��˟�ڇ#`c�E�	y���1De7`S�vr�+;�Kt�%k�.
�"Rg�&In�"�Iٺ��K��[#�Qd^.�'�Fb�<��f�d�M.�R>��䯘\��xF��B��W"���`�:E��������'�ğU�($�"�U�[��r��uv�V���_K=g�:\���vA�wo�>�PYh&"�%F������EB�N̷�|�e?�CY[�Q��}����{��]���X��/��Jj�(����8���7�`nؠC��Z�yx��O�\�5S�2�ǉ.~��Bcֱ����dO�soG��P�M����u9�ܬ�
k_WH����C+��YCzXr	E�_29�	�6sv���b��*��y��L՘`N�C����3�w����4��?�,)�6Qj�W���V@��B8%ڢ�)��g)޳ص��<(�m}�h�o���v�.�z�+@A'�6|S�LX���L��^\�Pݕ6�^��!6��YH���a`p}鼑��7������d��J���ʱm��
��Y�����
����H���oH��փ:��<2j�;S��f�nD�h/�i���Y��@�����J.S˂���1v%��E�kS+�QW@=�"���ղ����kB'[]��%8Z���'��=�\�z^����~��n�NJ����}�3狽�[H�u�g�o҄��o^b���7�{2~\M�p�젿�nM�Ƴ:��_�%��15d�$u�<��l�JZ����z�z�\�n����q��kJ���U��$���s� ��?k�<� ����E�8g&9lf\G�I&���0l���4=�"($=#y�B���-�E��>�Mg����z&�Y�i��u~VNCA���7������ �rc5&=Җu��J�k���˗峣r�����IQ�I�g����Wb���d����y�^ތ�v��i8+!��aV�F��ad��C��=7���2?
��%$�N>c���Q�`q �~�Z
գ�4�3]�|;�Om����#�Ǎ+�lNO��6�����	
�}��@I����.~7L!a0^	p(2@�%�K��gs��������a���8�Z�����:X~Ʉr.�[����mhsÞ���ӽ71��:C
�����Z�L�D�p��rC��n�6�(�����O�x=���i�e��_Z}��c.O�b�Zد����Z���Y	��]�_�/����VEz2��~ՈC���]vԌ�0J1�0��uv=�G���}�M�����&e�P/o+�h�P�YN%�O�0pk��AqW:	���}Y����ݯ�/�D.�#��=_�;�y�<K�uqʡ� @oG�	}J��kwZ�W���
E3o�{��q�0gDf�;L���~�Y�"
����!/l�'��E2��Oʅ�J��H�%��[@*jRs��|h�챮n��0ʺ`�ܔQ��[�qP����%T�y�Q����������|��]�u�%'El�ˉ��a�t��nzwh
Ԭ��f� >�DJh��a}I2ݚ(���y~"H��ʳ�W��A(�*���S��Cl`�5���;3�D�Y6`y�4k���W�ϕ1t�����`mQ��g����"��S%���qa2����G�Ё�d6��>m��'����P��4�M��m�ע=LW謟B��_�1#J� �"�B��s���f�Pħ�U���!Z�ҚL�TP<b�gc��?jh�=b��~߱��2�;"{	8���^���!����.�uT:~�}^]J�� >P*4��&dݜ�y��g���,֒����GJL��V(�kk��[��Q���L�>�`_S�4˂�V�,�f	��*��qbngE�G�`3��+Mg�����8%�ҁ�� 7�����o/�=��[ �5�b�i>5g��|.Q
�;J���'��z���=���ڛ�t0/j�韴�MR�M��7v7��]��_s�vJ�p��|6r`Ȑ�˫�qu�}�h��V#fǾ(`ͩ&�Wԡ�f�O�Ԑ�mi�N�)7���_0h��7G�M�\0��Z�y�[q^O�-�/�DO�N�7���,)J���$����$SD29Kڗ����#8mJ�)C��WM��T���}���ʌ�$:��6|g���وs�Z��p����)ĺ��(�����l��u��Q�<��>��$���::7_�;8�w�q��R>9�؄2L�S�#���0�����\�z�Z����T � �iHzhZ�L�@:*���Kfɣ���G����
,e:DO�9�ǻ�,o���+��Xs���?t}�v>/#�-wA�۽�_��)�d;]r�īG�7�����A"������^@�\e��h]�>�=+h7���������C)����^��p�� pν�f2w19�{ ! �-�� Of�����p������ĉ)�C�D����GH��<����"2O_K��_�7�?~�9(� ��C��0���O��7w�b���y����5r�@��r��Ct9r
�<(U=�,�r}�!-<t�cEr��)ӑ���l,�>V�/XPu��ȝ^�Os��-O��:G�b�v ��;�$�=T6�p����!u���0���:����:����ZT��}��8���~s ��t~|k�=�>��ݐr��d��;��ϧE��=GJj��lJ"ܺ0�i>���Z�."<*-N�� ˙l/���8=+��T5���Y�|��)�0ުÏ�j���8�h��3MĐKXrK1+�|�[���t|(�8�m7����_�>1��M+Br�����̡�*T�ٖD�d�M��4R��:7�<���3R#����&� h��P��F40`B��>��H�җ���%�}j5ֻpt��ȝ'9��O��مG��RD|���
ޤ�a�ͲQeh�������@<|�i�V֣L�%fr��|��	��
�Ms���C��ߎ�׈5��P�n�
�!ݯ�2x��g���J�`�����Ğ� ��ez��M�e�3�����ɜ����;�<{��o��L���R׹�>�{����턧��I%?c�`�{i�溮rv�k��T�{�b>H�1�d�pʇD��z��=5�:q&�ȧεs��/¦4�e��؃��z�(�&4���\�U�� �V`�����_#p6iT]�LӹT/W:��eAt�9�q�R�R`P���i��k/��(�,�TH��i�˯=)��lC����A�;m���i�ÕН��,�Uh�ߗJ�j�ڙ�x6�g��Rޥ5^R#f����) �ij?c�q�չh��{�Km�G��4J��ה3F���y��c2�T�\=��f��mW��c�l~h8ؚT"��[p[�]5y��Cp���b��#���#1�;���Ɋ0�(~)\�N�U���k3�,MG��!�+J���I���?/
����ý��5mQ^��X6'a���Hπ�KF�8���$�k�8)f��@"�͌7�f�[��*�'s ³ٿg� ������V5���O�j:���ϻ�q� ��"��9��Lp���ޅ�}B�R9/{�`��y�n$�����)W�͂&j?�A�W&��@�L"T#ʁ�ƺ��ĚS����~`쩥�fD6.��̣=�hs���N��d産O�ГW��/d1[ٕ	K���Swk}W��27�+1z-ҩɑ��34kǕ��; ^�]|��ɉ�V�V�z�
�/S�]��&�& *h�y�E0�r�z�+�qP�7���QĢh;��_^n�����7��!����8���.���Qz�b)�k���M���6�Թ'�V�'�(u����z]���8��M�(�#WjW�򥅣���ח#�s����CF�F	�� �T�������^u���+��h-}p2�+�qL\+$���l���;���0�w�����4�9̘I�dSfLw�!�5������<�sk=���#. <���nx��A�y�HH�c j� ��e	�U��6��C�Rg˄�fa�����f�n|�aq�E1e0�3�z���]��.a�zz��j��� ���ʾ�ٷ���k�B5y<���0�;c�CV����`��b�!����������7u��"�x�95�@��>b�_���@c}���ow
oǖ���������a�_��0�t�{f��n��E窖C�zk�d���#FP�ON����ې��c�p���_���T
�q3��m߷U�B��#��vX�+��j?��sT&�5KR�ߋ�����`�B"`#�p���tLC�^��gݍuK� �� �XWyk�m�]e&�]�V�:鄥9F���"Dtt�4�b���.T��(6^B��I>F�5&��	���v�����-2l0Z�9h�Uf0�34�NT�l�UH��M~:�'���#b��� 3_��|w�Ci��V�Cg�"ЌQ�!�d�}jZ�+0P>����-vZ��I�cC��D�Qۥ�-��������5�l,{�����y����O��l!���E$~r��Ȁ��x1��� !�H�F4@�6|�Ρ���y����}*w/��ZD6b���*��`����^Ǵ;�J[�}�Rۯ�ҹ���w����z3Dp��*�f�hh�h�RN�p�sx��mG�A�/�/�`~���p2�s�u�)2ƶ��C��[�#�p�QA�������BX$�#Wga��T	iK�:M���q�P!W��m1�F��|LM8s������.�J�!T���yL��V�	�kHK���Sz�U&O~��j�v�X!�#r7I!+u�������@�O�@�����-�XMV�c�D$U���۪/����T���������Ġ)��	P��3�-"�1������tn��i^ >Fq���Lz���9�O�P�ߝ�_�j���Ǻp$0�4�W���
3�g3��l�����zr�D��`�Y�S���}>��T�ʶ����"�y�*w�;ʔƵE2 kP�;���ݪyz^rܙ_�2�����dw={������{~s�	�<ܸ���c�G��v́��5;f�7ZUTS�A�?�>��׹����ȠoHE[�C���X��@8Xc5�5j�o��rV]�e܄|�m��&/6�J/����q#;quT��b�[����Y�F�ZE9��j�j�6��nO�:ɗVu-O۾"��Wjt]�FE>]�$�������Mէ�숰Fbß�x�lݨ�#�|���^`A�֮�:G����6Y�$�`���9ؔH�GgF�2-�Y5�3���ʴ�����a��N[B7�k�<�+K�.�aq�S�Y����s6�"v���X�CVT�����k�V4�%`�o���q�Nܬq.�p)tsu������K8��a��B�#ѓ4-�a�	IS���e͙u%2��������YO�&Z@���dd��Mv��oJg��u7�7��!�>��KQ�8������-�υ��z�(Ys�y��$^�y�3�d�����w�n��+���:���Q�2��:��_��y��pE,�&�����gW�`�r��ߓ�\{�G&�����sP�
g#�V����J�=�:�W�L��c���$J�m�GW��VS��۳gHU��xO�N��
�:�A5w�F<F)�eo�G�be%�h���C0��%r/�������)�g����/�%p�u��F��]��g��"���xE��w���R���:Đ�v�#�@�N�}���;��n9=?�F�܄V��VT��B�M�~kA�AW�߼O:��(e�$�O�4�h������]L���vu���6B�C�4F*"O��ϘP���.TU�0��W'/�3XEL�>¸
<�(�m�o>yw�d$8����Ӝy.��B��:�AI��B[�cg8p�1mX���2���DO��qC���F�'�X�@u3��{�vZ;�@����y"]�+��n��-���+"�ܯ���T"+�%�w?3�V�.S��R�u�����R�d�C���1��XֹEv�Kl"y���vxc-8e�]Ұ��W07�*�=���a�#���0��7'r�n~�ٴ6�o_���e�&���ܘ�f�,�k�)-v���z��	��5;3p5��	^m�yR���H����Df��J��JȲ�D�+���V�7?�n��^�n+�<=X:��Aiܚ�w�9����fy:�}�?W��y\ĩ)l"��ޒ����k���S�w�?�=��~�[(}��Q��XP��+,`5D�]�_f'�XYV�Ȏ~t^����KV
�OC�wdyv�E3v���9t�O]�`%��kW!n4��??-I�~�ZU��W�S1�E����0��^��ř�x��f�&��N��U��pV5���&ѿ��E��#m׭�&��'�6�q�(�L�h��O�	�@Q��Y�Epn�Zg��ڴf�tM:/�7bL���ͣqq�c���Jz���Ut�-ri�*F�1f����wtIx�b���?���
#\��s�}�k�M���Wi�MP�� 玬3������뀐ā3s1��ޑx�N��D�YT5qߓ#F��>�q��y�{�����lW�ga�wG"�g���ȁ�VҾx�j����`4d$��We�C�'X3@	���%v�1��C�*�Z����oΪ�QP�t�B+`y����N����|����
~������KƲrň B�r�9a4���7�l�xN���d�~|�F/��Y�(?F���6��ao\hUx:�<��Ú���j�B��nʨ{A�p���z~A�����������ȲZ\��w���5��K!2��):ҟw��p����`�T��Ԅ�>P�+�y$׍�$�;AB�t͐,�#&[$yc��Ki��0,���[�����ce��~��T������)iac�8���s�0�/=`=�:�o�����s�m	hd"u�ߡW���.)��7aIC^���p�6����w�XAy�,�ԣ��pP�Kܨ��:U�`'j�q�T%��ϓ�׹6�ZR`«WR�PLs<H��Ʋ[^n��� ����d���:���λ�k3D:�B�%gnet�a�����:֥��zJFm\����qn��k��
����Wm�G|��lJ�)���� �q��cPB��u:>�l[u(m*U���V�X�(z@y��-�ֹ�kQɘj*�����g�?�C >Z���_Ċ
�}�1�h���_�5W�I�ȉ#��	4�Q]��$D�I6���M �&Ϊ���1Yģ8���7�.�]VCv.P� ��X�r��0X# �{���!�M��t�� p�.����Nꯡ/��$���k�=��J?�*��߇�#���
P��V�GTJfw��ӷz�x^�O��R��#mQz<��/���P�΄w/���W|�u~���6@��W*���!�AX"X�i@��	��T�'���,�@HhW����W�ƻ���W���8<��9�Ӻ� �[$Au�?�ѹ;D���9v�)�8+k��T������
]���2��=lzNJR��
ѵ�yJ�߲��x�;����i ��ZC1���ˬ��d��X�8��U�Bĕ���PD�Q'�ה� =k6�eI���i��Њ %CaW�4�F���eJ�;����4���EW��	wɔ�����@��3c4(eF�b�����?z~�k�6^9j@���/�[�A��J��� -x�X�6�����k��b��-<��X����iJ�%s3Έ=x����uy{!���7���w]�3��'!7��&����_���dX��B��wx	v.1�T���'M�����iG,��@�[����\�����l�����o��d�K���fW���]�$��%��>�!� R��hYm��=�������S)G�u@��O�@:.��o��IQP	��X'�����M��'E84��:3� �}pȐE%�DF@�1ҿX��T���e7_��5\� �fK��%���zs��*�Si�f���L�}��Hwm��k�-e�9��Y󿐘sDk��|٪��Lc��Z4�D8Xlm��s0d��o)�y?X}�B���&�����U�
;�?"�R>�C�q�s�Rf�:�`�K9s5�����[���#����{�T�d�;\�����G�,��$4��sk���G�aYi:�h9�M�d-1�i]��s��Tqx��cP>��V��^7s�;IJ4XTs���"^��,4y=�ې��~�Zݰ(�����%P�������ۏ�t�ޞ�z0�Wj[8�8��"�,ys��f�>�:x���O�6a�gnbw@u���ೌOc�.Vo�w���v�� �ӟ�<5�;��_¿�0|�����d�=����q �%��<F�%�,M]�\81�������'eץpN��$��迉Y�u]�U�ZөY���n'���<ULm[|��<��(���cC�^:U��ID�%��f�e?�5�R��#��~{��t��T�����3����J�6Y`x�L%���p[,���t��z�2w(�)��7�H.?�K���}5��_��p >�*���Y�D(��U�V����\�"��Ŗ��L��!TJ��i�rpd����swZ[�����)F�$�f�2ˎ;`�+��򼳲oO���t�)�א�F�B����H�����$��p^d�dk���j��8k�wi��ppq�+Z�y�'��|�f���e8���	���`�˿䱣�ˇ�5h�g5x��˘/z�yΡP��<9�8�PnEY�B�oqM�AzS�ًQw.� �W[?	ڰ��`#}(CK˗��:\�D�AW�Kj	�[�rm���r+��q�c{'�^�?��3�pG�"&�:�ue�7w"0+t�Y�[�=`M%V�̊�8�����d?M�UF�4�cb	��;��2ϊj �R���!���#/�U� WVR�Y���os�z�wu�R|:��gZj�:`��-l(y�)�X��+�����!��!�S�fA�].k@������/��_�NZT���ޡhu�Bv�m,���i�i��N����>^�5�Ȅj���N�Ҽй"���aӔ!3{��Qg6������w�	��i�!R
K8(�gˎu	-3Mv��\�m�r"Q��ʲ|7�(���jUj��Q�S�I���~,QJ��,�-�|��9 �!��d�E�C��3�@�x���g��؞��ǐa��*��2�90��-1��Ȏ����Q!���*M�2*�fTy�i����|ye\�����T�˹�Z7�득a�Һ��A3�i��}3���ڀsa��z���d��O��$�O$��ģJ�ڻ�'?x|��Ҏo5��
dkafW�V�B� ��󫘒MB���-.kҌ*/��v%&�)7��4�Ƅ_V�/��F:�����T���S��}�(���6S��i0�����<P�E���W٥X�)B�Sn��fY���1��(Ż{&!�U��"��g�z�H_
����?&
"s�F�\��f���5�x}���]=�>_Z*��@�`ޜR����"f�RSy�O[;t��Z	�`	O�۞�<+S&߯��#~p9�
k��&�˸EF����FѲ��.e/V�r�Pٯ����\����=�X�X�Q�,>#J����\2�I�3����VJQ�73	)T������x��n��]�@&g�=�p�ԭ0z��넠��U�{U�p��3�?k%s�w�X	M �X�g�����C���OB�(Ǜ�C�cB�q� ���K}1-�Gg���gQm�?�4�BR��is`�r�������� 4��k��r���� )b�p��x����y�ن�F_�_K	�-�c���6��\0��~F����0�~�YI&���u�p�m��M��+�f�P&��Qd�X�^�wQ�j�u�{����˜w������,�k��X�}�J��K�Ӳ�fA��H�=.�v��V<�::7�g�y�v�el|��>���DA;gYB8��C�U�Xt�����
�W�Oz�xs�L�=g����!�iW���OX6�[�]7)Z\�dK|V⣺��"��݊C]���� �2Mv�K��Za�7�圌ߐ��)'��K�7H�����#�W��\s(-{g,Z��P<7`�(@;��A�7
�!Bi��6��!��˘�B결E��`~���E��]�[J�j�6�3��b;����`EF�n���;�nU���A�DN�k>��0J�B:1���*8s.��m�r��i����6���.ELW�+���!��z�����34�6���G�3^,�!�����8z��[����=�@Wk������F
pM���s��H8����/��5���;�	��a�v=$��#3˲��sP�r%�"�sJ��@�kEe����i���W�:(Dq�
����ʍ*-M	���>	������� ����nP1��T�1^�F�6g3�V�q|����ԋ�ۋf
�@���1����ϭ�.����L�Yy�r���:WԎ����I��5���.��!�ve���.9MvLpÆ�}������K�)$��6u�����v|b���>��vcA]�S���!)'���y{K�9�Ϥ"v�ゴד�K	�k�r^$�Plb ��=�>�?"���>T��t���7�,0V�������ܞ�q?�F/�b2���|�w�'K�P�S��-U�����f{4e�8J6*�ȸ��ͺ�|`��{������� �p�`�s���S�0���<vWg��怛bU�k3t|$�,�)k4���ZYvA�Vad�����^����[e)ts)�~��A�����N�CS���9_��D�`��;�O���
���LMnx:(��po	�����U ���e4b#�S�Vefj�[����P�,���M',��'a�ִ����Ra�%�OT�|մh1�,�ܒZO�O$�&Q�6�Z�&A�%���HR�ɁSR����H-7�g���_3
��s�y?
��b��V�
VWisU�� b&S5J�m�7��'�ۑ}ы��İ5�Pt�A�U7V|��9�?�%	b��(q�5!Z�Nj����V?b\�Ĕ��&�ZZ��:,���[^����и�d�hay,������lRez�B�ˡ��=�z�. �X�a�H�<ߨ��g�;����N��¶��z�M7�Z�u��W3��9QL$�/����[���0[�ry��m���;��D����܄b)]L}�r��(�M�<A9����w���yc'#����P�==Gp��0��r��!�7Z��#qSg������ߖ2ڜx�� ��'���(GT�����#꙰�oDA`�)3����cV۪���ȑ{֑Ύ�z�)�"��eY
M(��uB�2�b���f~�����,�����@�kG]�X�no\IL��Կd3U����� �x�_�6��gg�7:0#Hف�>,;��g��Z0��X���+�q��D�1sF����t0Nz��O�
#�����˓J6,]��~�}����i͛���¯��_�2\��W�U��	���,�wQo��#��!�s�q��s�c<:3N���I�&q�r�V̰d\�M,V�+��'&������vZ}�˖��f ���
Vx�" ���åb.�塔����h�Pi��Y��u\z� �<�Bܶ�0j�a�V�7�,9�{|-��X���Ԁ�(j�r�4Z��V��>dnO���%����3�m�Q6��+��!�D�Ip��S�
h$�v-	nd۝���2K�Gn�wL�m��~�E��x����ė�V��C׸�,!�@L��L�o&��=s��&��#��_`q�i��r	��w���|&n�zoaZ�b��$%��a	����u�y�h!C�7n�g[��֍�݁;���:G��,U���� ��[���م� z�hNxi��@|I��s���0VJ;V[3D��ռ)�kU�~�)k�Ne�?�8�!�x7 �j@��$6P�Q�P�Q��V�5�(9�.�Q
��ԉ��R�F�ٍ�"W��M+[���3ŷ���G�X�QB�9Va0�x�[d�ͧrT�L�!a���mV�gv D�Vy-�}+U����TO1�R@�*���s�D�G}���z��N���j�ˑ��8B���4AT���o)�R�\�^�l��?朗@q��}<!-�`�^O'|�g"y�n6,$6�rU���0dQ�U�ֻ#�����z��k�C�Ib��TCx'�Mrl@�y�9�^�4��=��0K!v@�}G\OZ�����SV�u�?����Vi��c7�O�3�����4v!����uk�߸k�K�T�; �ܤ^kt?��~���%��#q2�]���O\޸j�l/+�ռ8|�����`�4���Ï@$Q'���>��$�=��䗊T��RHe\�����CL������V
����G4j�P8"����Z�Ǘ��hg|��Զ׍�QEFc��6X4���t����o5������A�&���8�W�i�,[1�d�LB��$��t�4Wl%�iŻ#��2��+�ufI��_�*4���,p�"�1W��R�Q�[w���@?r�G��A�RNݗ>^��?Xd~u5��1r5|Ͳ�Ͳ�#5��U��vŲ�~�*��	lL5�����.�^8!r��}��AǬ��軤�T~_� ���ʆ�26�I��$���&u�+�M����qa�9 �7�tlw���f�Z&EéGDO�S�^G�}(�s�"�7�!���]ʎ�������F?��L�2�ӭ)�(��s<-�f:�c�-7����궴����a����L�\�l@I2�ŮO|��C�	�P���-g�A�=J�J���g���;r㘢���W�?T�f��ɕ4]H?����+��:��)N4��c���
KەqQ��e�h��s��-��/�Η~���o�5x{sB�ܙ��>�E�5i�eFKz����\Q�Z��3��S��`I������y1E�bS\l׭?
;���M��%���lkIth�u��L^�2<�T&Dn!����g���b�l8wO7K���gh����&{���h%���� B߿t���Ib�����(` �Dz�/�&|�b5j����S)/C<���*�u\~�W2���b�A'�	����Vr�������^��/�cFg-��T�@P<�%ϫt
\L�*��^�s_�`w��D�ov�p5�)@lm�٬!��P�{�I*Р�2���v/�=�r�7p��C�D���I��P�ޞL���]�������������DXa;��G�C�[�f\����Z@6T'XD�F7�C�O1b4����w}O9���+�Q��SU=A}�H�M�O���!��'���:�b�*O��4��Ga5L�SYy�b	%��+dlC���z�|�@��;�wDv�j����FI�.t��u��ՕNk�g5�~�5�-��C�ז2Y�Ȃ�}�`GZ}��U��?��G��;�Y�P隷ݨ�7�L��[n$>v���0̡�n.Xb�� �z-��)¨s�2@�f��E���M�S��\���<�{�+�*
� +R�q�w��b���qQ�&$�'T����Z����Q{����z�"jo�G�T5�nⱜ��#[�4��o� h�J���!�M��`(;�c��á$u��Jj��ચO1�dԏ^�(��y�����eJ��c��|>$'��l��P���s�'�q�Q���Kw�*�
��J�W�d��*��鐕�H[DO��vV�x�����@�`�7R=���(�S�1�GV"��T77�D�֊2T��%q�P��<c�y��V�U��� �,�,g�`����aR�>(G���s��R1KK���"���Y�wZ������Ȇ�>,[�@��F�%�Wv�ѳ�-ժ��H�ffΚ_r�K`HN�P��¤{A���*�̖o�>ݡ���=P�I����Y�\�7�L� '����v*��}���t�5O�_N����)�{�w2M�3v._�i*q�ɴ���!Uh�kľ~k���O�L΁,'*��%��Ԟ%7s��:j�j|Ф?gu_'���a�N¯��w�W�m��^4}٠��aֿCM� �]h�<�)S�6���7P� ���fZ���k���}e���f��PrJܻ��X*�h�n{+�_R�[��+x3o��C���V�L�~wvT��l`���#`왰d=�}�~�Hth!��a.^�O���x�a:.t�������I��Y� �H����`y���Ph*�(�����fCD�ޯh�e?�騟5r����	�3&o�.*�F���&첑�혛T &�	Ĺ%��ϙ��"�L�؎��J�j����ϑ8��uRt���[����3���c�+sj7���2!�e�R)XA!SQ=k�X8뫳Rff�UZ6�'��XUL>��e
R��w7�1�%�ؙ]QW�����q�Ax8����JTd����4V3{l>6����|wwD�q����������$4<�'&J|9ݖM�[���k5�8]�cvu���e�`�X�pGTfx$>�[֫�>}�m���3�w֜%��w�P��6��������jP {�3�'���.������;=!�ɏ_g����O)TYV^��`?�Q~:ubsP���
��B�o{�˥�k.n(�'Y���ʐ����q������
��.S��b8���EG�Jr���4�&(���ϡ�@�.1����aj\��m�^�ٙo�q�~�2��N):t�������6NT:���ċ�O�X�R�=�T�"ɐiq�e��i'#)��j���\{
��0�����8m�4÷6oX|¯)�3&�(��� �$R��:+$�˥Mߋ�	9��XB�vC�q粨�6YDs�5�<<��a�Cי-2>f��mO�A����@I���<hN=FA��o�`�i�3���2�ɵf2Xd8��\�"I�)x�)�u��e�g}a<~]mE"�O�ऐQU�y����3�,AY�S�=�G}�2�IPg�v"Vo�9 �<7K~�pFAa�Q�]�����N{7<:O���o��yά1Ǟ֛�BB?�D]����f�6���/��*e���J��0݄��f��_���M�Iͱ���j�(f_��K;���f"�	1C����;��G��[[\�m��j�J��q���� ʱ��0>��Kqg2/\�%���1q�_��0"����\�z��E~2$o�?���D���Y�)�.7���! �0�+�;"�]�S�.� @f���~���Ƽ���z�a���ė�O��	�W��={1Ҏu�2�!cՑ0��U�6h0�*k.�-���}K�y�Ć�e�sK���!A�9.,�3?���yD���?#NO�������d�rO
�����㢆7�,ݍ[�/�9-\=E#N:'���1�d�T�،��z�t\��p��š畢�.�*f��]�<�5�ɭ|���j?� b�Ǜ��u�죬����S��(�i@v���]+.Z� e�^��.r7W\z��A�sK�R
�R$qww�I�E�aA��3鈂��`X�%E�*�PT�����n} �i�#�fK��-��Q��36i����<�]~�1I������
�Cj;R�����e�����aB�Z�QXev����[�V ��O4z5�s�U��z��"��F8�$g�ʒ�Z��i��W lR��s4������T:]�ϖ��p����}��}�mxX|�ۣ�g	�
JXē'q�	���Z�v����!*ZX+��>j�ܑh��Z/"ͧ�L���zs���Ay���'F��L*��GH�χ<!�ǋ@�9��������`R�����Y�Vj�d2OU���E<�U�h�8�X�y枸 ����7�G޺����x&D1TZ���AT�{h��D� ��"�e{m�N���sI���6��Q�(X�y#)�A��a<PR��m*c�>�{w7�`[�ǒ���)6F�7:�qV}X>���?���Aw[��j�!V�J�z"��e�O*r�[}5T>�����/��!�Ī;?[����*ámF�c�bJ��������_p�2y�%}�s�Q���VpȾ��6�g.ɺ����*�	����a����c���4Tk�	�`�O�ơ�8�i"_H�ì/Ym�h��m��F�)��Wx�����}����BX�a�3�X����Ɛ�{���]��MSַn��p#XtmD��5[t�Z^'�l� ��>�>f�p��()��!���H���v;`�!��,ߔ�l����0s���b���p3�|�m�k ����jG�A��1��������R�7=B���5��?�i��%��N8�x1!�LU�Дw�P�o��\���E��48������>l_z���q,2����E14l��@H��u�2�C�`[�(m�ܤ�b�����%�3O+�C�E�hk��h	���'�ʎ�v�B�`��$5P���ĆB�p��(�����܁'k�����i� 9fK��ȌC�@��8gj�5���*aq��b;|��9,���R�E��I�K�0�>���7����=��<���c��X�޴eUi[`m�䭯*=���Fj�&�ďŅ���T���&Į�M^��d��ݲ���g"$�"���B]�U�;yB��Zj<Y���=K @���\ �T}`07*G�jԖ�!�v���9�\��D�9��J ���Py�\YK�Y�V1r�����(@�9����(�����,J���H�����ѣ���[l��'H:Qh�AGГ���kG��'"��p!)m-�G��7����h��c)����W����ןlO��/�ՙ�\����O"�(Ŷu�EA���J��@_H���	��ai��hE�^\�&0�ک�A��<��F���b�y�3Jv閉lo��^Ȋ:*���22�=<񡮭y5g��:`���}���3x���7��\k��m`9��Pd4�ExD5��x��+=��^��*�����!���M��R�Z ���9��;F�"��mz��m��]���� �Ν�<uu� \R�����񗺁���W:���7z-Rp�Q�	��ubB��M/���%�ɄE������=���@B+ʕ��GR���@�`ܮ�U���#���_b���O���}P_�XƧPD|�q���܊dbF�c[�g��H��V\����%�'W>��4�z^a�)�i>vY!䪁TL���?q�2Ũ��Hm��������H��KN/=>��ܴ�������%�do�e��BTJ�IZ���ҠS�sL�iT��tg�FO�{�9�F1.x����v��0�Sf�.`��{��c ��qE���+�6́o�ѭs�=\e��k����"c"mC	�46�fԫ��M�D��f�&�)A�H�Y%ي_��zZ�xvR�������:�):Y`l�p;-Y}v#y���{5�u؁�Մ� �g���<B�o`�*~��W��D��5A$�Q�F+^���b�=�\j�j��v�L|�艃kD��Ǫ�̥[��H��5�E "C��ZN[�O{���A}��2~��wo�GU67�g����xh�%��hRl/"��7���W�����4�p���?�o�Xr��n�_�$������Ɋ��8�`w��Z�ɘ�<ǰ�����6=������Z(�`�3R /%�K�0?�NT���f~w�M����7s.�F��t/=�������xT�f4n~��������ٞKy ?C�j��FoKIA��\W���	!4��>L�"�b�^��!}�鸔$���0�0
�/���t��
/D����"�F�Y,N�	����O��c�F�m2�����k��<?7MƦ�Ր�
-�� ��ş  P:h|I����L�؁8�P�N�
���H�o��d%J\05'c�������\�H	�Ɣ��~f��כU�g���5n�ᄅ�;�c�§�u�]c�24bz^~4P�N1�k4[xd���
�q�(r* �w���C+ø��xsQ7D����瞚o�>���E�'�q���ĤI���p�K���b\�1YԸG���sI���x�hdm��\�v&�pĽ��{+��kV����6ӷ��K���C�>�����B�/rU���ҩm6R���6y_�^R�A�6B�1>Op，��
Ǘ�ê�l�F4���?6]��c"��qm4wNl�׺"A"M	�H��j!��`y��x���i)�"U�lz�i�l��W/M�vUlX�:���U��d�Ct���!���-]uԔ�3$�F�m�{q�>]���i�Q�\Ŏ�z)�B5���~�а��{��P
���.�X���Ⳉ�*4e���G�.3��(f���Y��Aq����t.FQ�:�x�Ԃ3W�>ks���
��v�͐�W&�j�Ct��С�Ug���C^}���4*�
�J��xB�#�g�{�j�	� W\E���|5����P�p~�$��@������%$�4�^x)~�oR�j�@�2�$o���*X���^4�L�����\{�<�2
�~}ffL&�T�Kp5��z��8��B2Z��P)���bEL�>�t�֪�ޛ���nT�l+��-�#`k�Y28��J�@Gg�޿�1�d��(�$m3	�뺰�k2ä���n���� 4�������8�خ7.�}�KN�˔?��
tB�-y��//����x����۬�^�Q���4������6u��[F�zh�1}��R��c^�*��-�]rT'�LVq�	}BY�Z��N�n���OWֿ,�Lm��=�0Q�ɶ'*S�W9!�}e�h[�*���A�m��/7��5o��j����'�֪n��#O2E��N�%�ר��$�URl��o��Й���n]�o��Jy�+W��� 
\��R��^U��X� <k�T�����J ?,���iTڹwˇY%�����%qv(����LF/�Ԕd�΅�c��#�J����y��� 2@+_w%�34
M%�=}mX��v"���������vk�B��/�9V�"��J���<c�3��6���18}A,�9�E`y�63�i��^�F�
O�~�m%d�5N3~�}��-��
��N{�%IZ'o(�[����z	Q�j˷��.�ͫ#��^��4]��qZi(A�v�ڥ����#$K������[U�4Pu�v_*D4[6�|vC`P�֕=4���r .���V5��`})%�T
�*"��)�|���%/2��8�ު:�m^���eH{gKK���!�f�c��[{�$k���Ƃ_ǏB�M�LV���9W�^�*.	��F��a����#�~lH�2n��E,����t������f���ߗ�Ꙇn��w�8=g-�Q��x:�O���ٰ������L�S��4o�Z���q�x��A�]�2Y�Ě|u���t�/6D)�.U\[,x���֔~�R��:���iI(�<�����*����5,A)�oV�ĺz7^!�W�n�ul�`\x�4���{+����h[�s��vM�|�B><�(毩��:j�jѨ !,���wi���>�-eևw�w��}��0��W��y��f,���n��b�q�V��O<�}��b�|0�#J/`J���'B�_�s�����c�̡���\Zt5���#LD��8qp�ɔ�s����"����m�c�|����m~M�q���t9��O����������`F=����tSv��y�'M�l��IzeO�$�~G���e-�1�����S�G��tf�����R�2�h�7b+�З;�|��0�]�4NWģg9��w1�ycRj$D���!0=�?q�S�/�ܨ�]���n��h��"�� �<L��H��ؔ��QE/���Q)��F�FJ���ć����N�*q.��ź�	S���MJ�to�Y�s�Jo���@G����Y���l���Аʧҙ��Q� ��*��
�<���5��Q�����D�x	�+�@�B+N ��w�*լ|����Kٽ���?�w�t���ݱ�|*=;�����u�����/��4�<#րU�Ne��FAʟ]V�ԵZ6��#�0 x�^�\�4K@P��e{A�x�%ѕ!�ڌ�	`��A��k/o��z�ۙ���V�jdԲ=�y+݂���q5&��}�(\�LX��F�q�kG������G/	��쎖��'	�:^�ђz9ab����iy��Z���	x�_fʤ#b��1C�����
�����CX+o����|����j�rØ�C5�z��N5HH@<�JY{+s�[fQ �Fr��E���{B�Q�d��j�!��R0p�49�W��Q���Yc�%�EirJ����Hf�h>��p)|�v+j�y��KcY����Ձ1���MY�����Ɩ%�Ƞ]�$J۴x�I�����<��I�J�F��HUߟ{+r651��F�x��fq�zϘ!9��P�D^�7����^��Ji�=Ɋ�/#���+���,zcnî��<�ݟIN˽�guJ�����=g�U�;:������8˕%�qU�킉�#�$��dgi(�+F����"6��U]l���WM��i(C�"w�y�	ȸ�Dd�~U�������>	�u@��ſlGM�R��g�yl���g�V2�cCR�����T,	ћ�~`u�o�#�ݯM��aD���ٗ2>4�(<�H�f�n0s1b���A�\����[X��{�;(��js!	W��è&Y�K9 �������9;ښF��� ���k�u%~�[p�M��M$կ�'g��9+գ��zj8/1�����x��L�U�pRn�:=/_pk���a";������@�
B��X�
G�'-- -���
��˱�i�{KJ�k) �n"�r�9���.yb�`�:]]��ǦiW��ȫw�B7�1L�I��Wr' �ڂ"����^)6�n%c�G�$[:$�L���t����X}S�����n*��aӞ���)ҥF�B�?�8��V�֚��V*�~�@����c���I
O��3�qG7��O�I<J@�i6%�/�t+t���Dj�&�\�B��Q0Zn���%p�f��h9�IMkC����+�$ �mF\�⒘Pȧ�2����x�1:{��3���1�Ŋ�͞z �s�LƵ�KA����.c"�t�Ɏ�1����C1<�K�?��@��@�=ݱ��-q矦�(w�?|3�j2�;�C�]�f,kK�=��r�vLĆfva�4i].���z��̒@�l�EHqR݅`G�a@�p��iq���q��o���Q��=ޞ*��p���t���C� �(]칕����Q]��;C[*5.���j�K�$�����ڜOn�LdW3a�`���4������x�\�p�?8[�X�����"�<K�)��@��ytqZZ�-NP��i��oX����~3�R�1M��H���n�s�<{�Hn���O�S�D��r	=�$V�w��Rb�'���ZF!,e�{���$�Z%��1q5�ر�=wz�,��ԉ��h�����/�)�	������%.�u_�ݻ3��$"��7���1	�o��{Œ	�m�:;.U	��ԫ��H�E)��[�Q�ʷ�`A�M�3�7�ƀݗ^�Sr˺b�~~��#�l+ʽ2�;Y����3��Y�t������8��h�e���s��4���?/�q� t�NZ�x�<�dBJ�}�O	�������o��L��dުk���w[՘��p�")?25�^�C��;2n���'W�Q�u?��Iu�PP5��b�ȡ��G�J+����I��б]�t;�m��4`��ŵY����Lӵ���,���@�*E�fޗa>Y�meW/�ܿx�ة5��c�'!��s�1�Ĉ屽�0?�Nۄ=�3�y���m��aN�{�'��Jnۄ�z_�S��3�`�b�������n	�%7�^�҈b���b����'H�G|(������\����^���w�>8���+���c ���'Ĩׄ6mn4��,���h#�,�qB�|�V�f�V\H��|�׭K�>�.B)v+(V}����Y]&�t_���h��>Sn0�wY_)^�f�Zx��n�N~��Z}}�%!:���}��Gڕψ�3џnNLY��.q�𜕎:S�
��,����ِ�����0%1��s֮s��"BB�Z;٧q��K�k�Q`pu/�n�iB���a�FP�~D�f���f�D{����]T)��c$I�w߄���u�?%��k?���g�����!M�����6�"m)��H�U�x�o�7��9٭������VX�PP�3W76��p�����&s���`7G�-Y:����)JX�c��#<F3�W˳q�P�;�����G��gj�' ��f6�M�:�]�3�Cnct�T.�9*vTu�=�{|&|��:#��
�v�Gq_[ɍsl�O: �Q�Sܻ�P�4�I\N����`U����(�����V���&z��'(�}�:��'KŪAG��r.O�f!|��[�^��4�o!���H��Gw�ߜ�	�2���#��B߷{����q��Zug�`(9&O*�$���+/֑oX������I)���ik`�/[-Vj�ʖ5���q˔�=F��ȫ}��h$+���i$���Pu�~8::Îl�^�׍9�9�S����6J�$��AކL���&�j9-`	��1���[�۪+�U�ˬ��~��GÛŤ8Mf��|�� �t^_�9L����}*��'���",_Z�;����C q�j���Ċ��4�TH�1�!��|]q�qx�a��گE�X!ۋG���7g.^4GJYe�m��;j�* E���eB�ctJ'%�VBWTH���i�������f�9���(M*�0#&��	-$ԭ<�uYg:?B"��J���șvq�P��[5fB������us�0�@�r��p�/V�E$����璨ҤKR���l��2�0�S>нqM��u���As�m�Q��8mv`&�?8Y��#�iW��W�j�N�I΄V����[��Y¯�g~W+��/�q�($G@Ґ�jzn]���t���VW���e�d֍������|�:ÆRH.���{��W�T��ߜ�	i���(h����~��㿑���'y��KQ���3����ك5ń�D6A�[�{���B>��_���	�����Ȏ;c(7�_���X�ߟф�<ϒ����ce�b~�v�b�)~�v��b�����pe���^��&�A��%�cG������^���G/��Q�۲rt��EE��_�d{^1ϐ����Ro;u�y�>�J���a�
��b��c9׼��ƃ\�  �]-������⡫F<=2���:�&䫉�g����Keg<(����&�`�?9^\�U�A�c�Z�� ؂�}L?O�d).x��2��߄͊"e_z��(?�G6n�Y��2���5rbՠPb�Dl���y��~%��)�6N-�<��F	_May �c�څӸ{3�+ya=G���h��v�b�Sԣ���l�����������rz[���9�{\�t�ʬ�����6��s�^�1P�N嫝`W��<�\Hw]���6����w�Z�nG�_�a��5]Ԑ���Ĩ��˽�ɟ�<�8���۷m��P���~�+>��g;��L�+�����<aR�G�;���	��-����9�C.�G̬�T��[Z׽ya��͒++)p.�X�x?!�+Y�C���ދ�]څ�C��N'�6���o��`��n�W��GE[�1�7o�>ȖO�'�THpG�ω�P��nq ����E{ ��(���hS'ՙ�@6�JJr�i�eݥ9�f���w�#v�1	�-�+���5S�g�Vi�I}��'�ܷ� ��n���5c��t��PEb �N�8_����]��������M�5���T�ڗ�r���l^�"�*|ƒ�����nZTO_
N��?�����,�~��PC�f��\f��H�w1T��3���"ȭ+~S/�r�8&*>�}ֱY����1�1�ʤ�~��C��gօ�@�Y/���\l��%2�в���BC���s�&��+���?���K��\���b�/y`1��u�5k�:��7v�Ԫ����֪�3��.�� �1Li�N�q9 ���Fq��p��/�3ܞ�a6�oއ��7�A�R�1��N��\��M\�Zĉ�'3.}L������(£<(m�Q���*ʠ�`k?hC���S�C(�u��9җ>!����b��>�(f2�G��'q����������T&Z'n��4%@���y��U5r#/2�Fr*z��43,ϋ�zE�;DA���%�L����n���陼��Xu^���S�(�vm���3^c�mؿ�у#e���� ��~$ir�rP��!h�����QB�� bJt�V�:��i����.\�2�[�s�{�&]Bӷ���V|�)��*�J�
I�t����&zP� cZ��.��Ȉ�P�O� ΃���I(l�N�@H%��K�)���$ԍ��'-�D��c��Y�D�K�IK�DLQ6/��e����pV�AI'0��)#�Q�P���#Q
���i�{���}��b���KEpX\ř�$��Q�G5r&�fpq)f*4;F�/�iR��>x�C�xAR_a��i8W�}&&:;�po"���lFm�����so�`�`�����e��E.�|�L��#�q�l��5l�J�R:��I,\C��V~-�=�s�]�c�I��El/A&.����Ԕ�D�#<@�7W�k;O�6�ݑ����rߑ��wT�}�VE�}M.���6�X|g��r�mj�LL����%c�m�ld?��SR�=� �VtJ��p$A��@����!\N�爛�|l�2,��$ID� E�.�E�pM�_���'�͡�L�QE2�fK�B�H����!	�f�Q��.�ʞٕ%p����zyU����m���T�פ���(�E����ʶU���{@�K�x������:��#�`{����b���l�8��Q\%%,�������
i��A�6dmW>� ��K�"=Ε\;Nm2d��j��KX��gG4�"#
f���
�t�i��-�8�[R�����I�Ct|�^ƍ��ٌ��m�mn��8Hm�_a�1h��Fr',���=gh/�ڪ/�����Ř��֞{]���c�T��}�Q;,j�z�M�t�ZGAH���oy>�ϠR�]ű�^L��
��4�?�g�F�⮪��9�k9�hk3��S3���{�
�S��l����v�ZPR��>o�-�ÀuF_�6T&C��Lj�#+����.���*�N����ǀ-^���8.�_������ДK��C@�c�E/���e�����I<�eF[tC3 �)�`�wZ���'P*��1���.2�7EK�{վB��c?;E9m6hTK�3T
��_s��s��n��S��#\%�M�U��*6.�/��"ls~��/�JJ@�10{�x�����Q�����L�]'7�悼0������3�cZ� ʨ�i�k��n����=�ZM��ncKx�P_@�fP�	J�����g��WD~A{�hs7���}��$#�Щ1�\2ܳX
����n�ï�#�G�N:�k�A���W��7̺�c��2��@�m|�׸nK�%_ymdCh4P��dr2���X)w�c7��6Ο��>ن���cҪ��@o��H;�6cJ�{���ŵ���=A�#J�''i�J��O:� 
'k�wʏw������U������ᲠR=��4��W�Hv:�^����k&{0�|�zGwLD�ѫ`���HG�l^/^?-ӊ�+��zm0֒4PP�|���_��VhL��H2��N�sfC�(���rT��dp�9�=?�#�K&� ��n�F��җ�OIF˗�;(W8�()������ipU_����.5ƹ���'���ե`ʳq�{����a3�5.�eE�P����j��Vd�I-�`ε�:Z\�6����3��� �2Vw���*��W�ڏ�%�o1�u~�zѰ�4ÃI�R��T���^AH��b��ws���NV9K5{�������?W�SlC]��mŃ� >ܖI�چF�Yl1�e�q�S��a�'d�Z��,O��Zh��U�� ȕ�H�Q*��=-�XrE �^Xq�z�}�0XH�.���h��Ђ��H���OK�_�%9�o,Az�*[�r\����uE9�����r�K+�x�R�2���;�Z��-V�8�5�
�M�; 2{����{fa���2�����0׎�����B�B��Wq��9q��2��iI���Y�Q:Ap�;�?W�p����I�F�R�I���LNLAā��y�w����W��h�X��P?�f��D�hd����+�8Y�ZG,m�^�[&1��i�v���:Y5�L�!�����ׅ
��<`�D����� �).���6��k*!.���g��Ԩ%�@�:�v��#� �ϒzdW� �]y�p��0n^�t��x],)ǰ�v55=���~�h��VYW�͔���7�H�e9�k�]���V��V���Ei��E��2*�J��;9)!���@x*�^D(Ф�`�@4��#;W9b�����3՘;��A�͠Tf�E����":��Uj^n�eK�8M����5P9^#�:��( M��V����Zf�����5����k����5���_�Ф�����y�o�l<�+�sɹ6�5AN��1���%�v�����{�7=���_��ؖK���\19�v̆$'����#x�i���#�����2�5��X�pLJ�t��u����M�7U���AKN!ݣ�n�vB�9܋H,�P��E��v��\E�"���Ӂ�u��5��$&b$L���&~���ã�-��c���a8��$����k�����0�!1��$�bR�nȔb�����	��K��F"��z������%�q[)s������)�jZ�i�a�L��`ً��=�\lب��؈�<��ǅ�Y�@kL�Fz7B6@+�|����[��}�	�����l6B��(�@���u���]�Y���m��9�=�:���K��SN{5c������1@AT��&�Y�-e��~򫻠X����,��#�X���_�ڰ,�����j���� �9�}V��iE��h�� \?7�C�669p��,�z�<x��h�X�|t�s
�ޥ��B8ܧT�g���*%�|),Uq6Mͷ>�Wzq��&�;eJ>��L�KjW�`�$�����}���c=�>@�<l�:�IL�����D�"�j3eU���.�����k�؂En]�"��<��f�4\��*�E'��f�}��v7���1�M9׮��$� �RZ[s���h��4t�����*o����u=�a,��{�\�[��nt(ys��"'I��f9=_DL�N<p���,�6+,�X�P~��I��Rd���7���ʺ�Ȭ�N�x���L�AM0mq��h�V�Ɯf}��ߎ<^;�}GS��.\�(�d.��ɇ��H��N��5� �8�A ՘�M� ���4>6��wdԨ�TG���+�W>��M����h葸���$U�L)�LkP��"$a�vQF�7;t^|�jJ�f^D���K���L49��3rBj��YR)�����L��T��������p��e�阾5�^��4����65{�������T�ݴ�<�X�KWJ��NI.:4�Φ
�
�?�8��Q}�;L�Jv	���&6h����~#BTv~�>�R��6���H��@9�(�[f����8"�nES!:���)h[�	�٪�P�N�\�@�ɧᰏ{�Sd�F�/E��sh�����$y���C�cΖ��	4.�/���*���e�	�~�0ԥ#}�5{���:�C�8���2��ٓL�-_d��i=%<��f~O�b�6�o��I[E�2� ���y��,��ջ�۠�ns'��{�h/��
a=a	32��ˤ�������}D��+��q����D�bw�ҙ�@:�e�k�f��&7�^���ڲ\��o���`AY���Tm�>��kc���
Ȼp��u� �z�t�ԫt�O�dV;
 j���Z����-�n�|}��"Ą�G�V\�ܗO!^���3l�������5 b���P��r���~�q\��7�T��u����c�p�RJ�Lکx������׷x~����������:o%_o�������OS�z�.��&�9G�#�V2�	9��S ����7B�B�&����=� ��Ǚ):��N�����F���io�a`�Mx�!�Z��M��!��Tl�B���̱�(���1�=w������4�N�Ϊ�o<	�m	1,�u��!�62����IbQ�`��Jbox&R��Y6/��Č���>�<Zpob<ѵpM��<�my�j0�q|����o��W@*��'O$$��RG��ˋ��,�vf܎,|�L��#��p̹�Tp`q��6y�U	�_�3��:�Z����SH@7�%���e麵o8�u����z��fU|�(�фl�>V��������9�ȧ#&+Sɭ�p�x˴k!�Q���3�c^�)�=�^ �fOuQJ]�F糜�\��9Vt	���N��w)��\�d��&k%Ȱ� �]O�Q"?&��C��'T�hym��A�]��3\�R�z�~�C��|H�`�ʢa͔�m�"!HL�Uo���H��e�n��|�3���l�և���US^�1��	9 � ��HPs
���V��#�B�)��2Dִ�>zV�&���t*U��Լ6��1ѱLY#xi�ɏ�,��*:�NoS�����dA��q�M46��%�D�%�V��� K�,O�ؓ,��$���1��X{- ��jG�p�S����'�q���3�4�EK6����a˫���-ӎ���I��koiD�WF�n�h\�j�+��u� ���N��w�d�@fjXޕut�#�S1p��{Pٚ�jЛ_(垛�̺���Ľ>������l�|2�+�GD��ו�+��2Պ��IF���GT (lEp6�'��θ��>(h��&A	M���	��m�3�VYg9�p�Ͻ���,�W�Z����O�������A�Ov�|F����*��BP�;p�~2Z�{F/��Y'
}��/��ǚM��ۑߗ䒅C�_�zWE-FmPX$,�)w����0� �W�ZR�S�S�*j�f�TGFe�8�;�9T,D��6�DMf=���c�"��Ukc�m�f�Z�v��k��q�>��Pk�H�o��HD�y_r���g�}H�2�/:qS�z=�)�F#c��U/^��N�#v���5(��o'�Yr��S��trt��VC�z���B���`�Eo� ;#y"D�xvw�F3�0�����b�[�@��n��2��)o �����.��p@�|�E�1�����Z`�B$ɂ���y}R��Z�$�u��,��-��y�����ys/L���R
�t��3�S�e��4������N^ӹ7�)D�	����/��p�8�?^��\a�Tƅ �c$䲰��LWc��][|�Lr�O��fI{]	C^��B5�������I����1�����Jgg�X�oO�l�uv���"��Xxz����V��K�?�	�'mT��J��C�yJvе���6wt�wd���<�b��1��*�4�c,u�i�g�qrp>��@8+�Ɗ�ĸ}�wN��Ŵ�<�s�b�'VmTv���h�:c�#��{������T��{����*>__cE9Ћ)�I��?q��R*z�6A	;�̏<��.U���PQ���I8�O^��&+��Q�f���7��"?Y49��8�|�J��z-����03=k`�Ch�%�:.�b�W�Z� ��{��D��(�����8��D�����q��p�ƀ�)�VE��9[��`n<W`bM�[l����)�ް�o��o��O
h���N�ɺ��CEg�j* G%e�k�$����������J9F��Ku�v;�&�PA�PM3���-��↧-������:6���-����9���G�Y�V*�Im<�@�`��\��9�"�,fRsP�cϒ��R�lg��P'���4���2/�?	_���������aY�յ<'�z�/��U=<Z����\��pJx%[��4K���z�j��8�[=�6&�g���H����w�p�� �9<��#'$����?��lU��UO��EqϷz���y\Z���a�Qb������U��`�|;�W�^�#E�L���;��_5�W{89�tc��&����<v���ǵ0���2 �<��41��G$����H�>n��lF�VZ]ѐ	��[�K�/�W�`�2(�(ˁ���ݔU$�ĜԹ��/�K�L(0a�_kLe �9��#c�u��B�X8vN����H�7a@vݪ��~���H��Y~���E9�����9p���'��N�_���j�<�������lCp7��;��hPzH^oB�%�()���3XԈ�HoY���)Xc�2�s*�&�*�>P:�။xu�œ�i��>L�΋����$z�M�ؤ�]�[�7�F�(�N�ɐ���`oM�3^�_�S=�s8p����I��!q�
��6,\��9���$�E����K#t��u�ȍ)3$��g(�	�ׂ� ���7��B����*��3'۷ri���?RƠ�ܖ��J锑���2ȶ����'H:fNx��|��R���vh1B�m�j���g�cZ�;ԙc��C��o���<��#J �>���z-ʷ"Rpl�[��+��f�EC��M��$��4l��M�S$|��֨�]D���_m��z�T��>�����H����]�1R\�T��A%r ���	�ެ����VR�S�:�K���`Uzw���r<��y4҆~��۲�γ�"�^8h�Ԓ�S ΐ�X	�ܨY;�'(6#� ���|T�}�y<W(�6���g�µ�	^~��5�����6`�Pr�@C\�����H͕b�"�[0���)	zݡ�fO�v�5 ��~>��+�quj��¦���S��Ze\p��7���ƀ���	��"Jϲ3��5��/�����5椶���/�q�!")7�q{�Ya?���z.~�ۂ�Y}���l�2���Xt��?%��(hF��n=)޻>���K�;�;|���Ç����T�o5���Ǳ�C]�Ο�cq�^@k�=�R�24�h;X�'&W��Z���/㸔�f'������4;�𷄱�����t��~��P�l���,��N kPgѾ�G,�ca�&<t��G���0�%ikŖ��7�u(�����(���j�=R7�t���y��cT�f��}�j&T���p���vEe9��)����mت�2�UZ'ډ�ټ^BΊ���ŚU�I{��F�R���9br��Yuޮ����P�˴�%N �a�p����r��(:���tE��î�=�ZZ77)�g�t���[|g��P�$�k���Tn%_����{߁x���^Mn�	.9����E�:3�Ot1�Kz��D�9g ��h!�F���K"\��E"*MD`�2=[B�,^�a%ѓ�� �b�����%�i��Nܰ�f����>?!7��Ke̇X�ԯ[�h��l�-�,]O��!HN���RB`�Qt�0���m��wp%$Q�RF��H(y�:��9a�a·�2p=�`UM� 	^��6������V�;��8�V���x��0����/b�2i �E�S���2�+�1=��3��_Q[ӿC�?�>�s���Z�!���vk��r���)�f*��T���:��ܓ"�E�\p�hM��ϖȸ��j+���7t�!����B���.�1��K_�ξS���&3 Z�Ȣ&@{4C>�8����zlCj�2�˲?X�p�����%�"X�q��K/�.��_N�?\�T��O
�!Y.LOH$z{e%k�`�1f�)�p.�g!APW����A��3.��iу0�>�{��]B����}6�G�i�t�B���'�R���Su�=����N�X��߶��ѩ8l�X���Iޱn����7���U��}�{��^]mi)M�c�^���յ��Œi�*G��'�JRN�LE�!�0!����?G�����QB���"y�c�r�Q��>��mՀP�\u0�9�'��0.֬ɇo2�BB��	�7��1� ���������ܙ&�X4���R��r�{�Ԑ(ڦ��av�y�W֛�6SQ���U�I`��>���X�\�#�&¢��f��d�OU�X*��v)�G��<{�~k��rKA�̥֬�Aȵ�������4xc�Ft��kP� ������h�Us�H�1��\l?E
�%j~z��E���R~�N�D�H�j(�k&Y���Pz{�ƈs�3�+�C��n�w�V4L�������b�۴�����*34��
��:�#�3�[�r�5+�Bcu$�������*F��&��泌�i&�QZ���)�3��şӸו�Ѳ����E����m���eqY�<!�'_zx�VZ���fǐ+�W�>g���no�6��c��L>��Ld�*��j�Vb	�x�x��Oi�l#uWm��@��W6H�E��M+����ͺ��-R����-������������ګ��x�h�J�3ς��A�4�"t�w�&V�^z��k����:
*)a����g~�������.���?�6�~��&�R/���CT�$��^hYvI�P�����ͳA19>p�*��"��9>�u��[�.Iq��T|�|��:zm�}��A�"����'�ɮ��0��FSmYJ�B�ZX����]��h=����0�2ȭzqqܼō���@�Z����'6������}�4��f���'&^���*�����r���	��\��x�"w���5ӷ-��Ӥ��C�[�m�9�~��U�����g�Z����J� �s�y�D�M9�
!Oe�m��"�s��z�]�z29�B*%��K�d��^�J��e�_Vzk�j�>.2}�V�?Ԭ:�~���3S��q�+���7��$�'Zh�a�|�H�|<x���g�R��H<��0̃X�)x�DΝl�:�,�7��5�|o�k[����~)3�f�k�/��B/c�uDC[����s�cMF?i�F�����c"ME�I/�k퀒*��\ufx��D�<X����zE��d��G%�%)����6���4�t'� �`xE>�;��(502L��j��s���Y�����+-1ΡF�+��?�\�x���GX����
�?r6���(�-�u�h�x���+i}�`*\�W0��P/����zWz\�z��~A�|���~8��z�ܕ�������)j
�������8g�\{���^�;q�[h�éSOS<�MݭMt�+��r������gN�Y�s�N |<�`��ڜ��M�a(ڴ"��}��π��#�q�	tB�$�i�-sA&7O.�἟�_���%ג���v 0ak��$w� *^��Y����@��f��6�i��n��b/�8or[����ϜJ�����#�N=�b$k�>/d�D7eYI�}8�c��:U"������c�,@�tQx��0���� 
�!��E�ځ��%k��o�g>�#M.S�F�Ks;�v6o���D9�Nҡ#�\�v�����{��p)?TFu��:�فF��-ɑ_��~�Gj���dy���Ҹ���mC��5�7����{�2;3����\�-��3vXӈQ��)~O��V�]!,UY�<��?b)���XF|�M����#��~�;2Ѡ��*wz�/��	�2���	�0@��x���}������(�z}�<&X2�򴅴w�<|�+�  4,����x$�j��gĖw�z����E�*f T}��u� �P	�k|���&?g�w(���r�l#4�tÛxwK���!=�Zi'51M1w��z�R���Hh''��}٬D���Ү�9�E��0^�Uw�U�r�n�&�G��h��F�V��R�U~P垡|��C1w�4ap�vu���g=&����ݫ��p��[�j��@i��O�s�°Z�-��NP��vҩЗQH��@x�+F}U��ک B���N��;p�ư�%���͑�|v͔�D���4�p��}ěc��T��RX<2]QD��r�d�������FV���b�2���"R��էN�e�z��V��������>�NC�s1�>�d�g�Ӡ�j�Ҍ�|V,�Q%���\
�A����4u���1�H���	��{��=��b@�X�<�y$,D�o�׈��I+�@+�]4%�M�<���t��b��5���6����Q���g��c�*�9ZIH$k�n�e�B�Xy8���S�+Î��hl�A�n�|�"H��R.����������	��n#�ƉTU�h;F�[��E�\O�����g���q r$Y^��g����""~��o���m�\j�$J��Z^R2%�EG����Q�v����\�K���6�T���]������H��Պ�W���������ãT��1�������.'�� py(�i������udSR}5+��M�-��}�TSogB�yĿ�2�HZ�ڱ�Ĉ���H���(q� �IS�_mr��O4���>ȷP�Q�v��/��?ө3`�b��n�����_�ݷ�vV�*.�v�12M���<4�S�$��v�MO�j��1?��RA��9��~T�{��CY�
ǚ1����fU�>T�k&�nJZ�>�)�
�~�4�r������8tR~��ӻ��c�'�=n��P1�54�2*c�� ��E������,3!J���b6�ē�Ə�V:5m#&0�����i�J(�5�����Nߥ���$�5B�S��y�d��ϙ�b{���pe�0�Z4�]9F�қ!���|ѥh]/?��������;�����=�+wӝ��a}�����Q�%����	'-=���O�:��l�'�G����[�}@�YW��+H�x��4���mM��p�j��v�<�j<��g��_���R�a�X̼���ﶪp/�̐yl=��u�I����G�b��Y��V\](�����e<�X"�tW�y!}G�����|��Z�|��%�И��p }�ۅa�q��.�>DX ޔ("I8�&�({���� e�R}����'��1Xw�(\�pD�]C�=�S��G@]�躟"^H�J�}H6�x�5O���~lv�OQ_"(��S����P|��6|��>+.�,cD.r�2,O��@?fG������#˚�|݇w����FCr�0�l�BSH�)h;\4��~�f���Y�w��=v��p�8М'8ȫ�����@�}�^/{l�N�tz�kn��������!V��T��fuIKw���N<���̳Pw�p�y�)����D�~��t�{��5���IQ^��JF h6V�yD�}0?-{!fZ9���4l�J�]WxQ/2�`��a�.c�Hh?5��Z�/� M���b�	���L%�XN.?���(��<C%$�'�38	����ÿ@�؟�$�1y�h�QXq��`����:��=!`
|�����4��p�,���������
f���Ś��hB^�`m�}K��	�3�Cc}��5�&����JʁE�y�=<���?��ϕ*�@�w�Pۢ���W�{ؒx�����Ȃu�H�c �ܟ"/��KB�¼vbj��_��8�@�Ǚ����Rj ��ߋ��K�E W��E���}(�G� ���7ۋ�9�c.,O~��t�E�������['�}0�9͇:^$��p3�'|bƅ��{y
]A�_��th�܋�����䢇�&���[N�y"�4;u���١&��P)����Xp���;�NuE87�ԋ)�Ł��OͦK���Ymz�֯r���K=�y�ђ� o�@�"�
wD����*Zc�M��/�⠳�N�t9�l۝n�:m{��/
�H�R���N������lͫ{�}��ey��{��@����9�́�5 ���o����A����jz��*KGL�c�qY��A�^�c�Ʈ�bLю��V�n"Dթz�y�u&���n ��xT"(�(��P��R�M����D�0��w����Θ������_��ɚ�8A���0��n����8��v���>��N��X���<D|��D�Ef�]t�A���������jZ��3�"V'.��c�3:������9�p�_��bE[,��΄y�)f5�w�3Ma���"� �]a�L��m`A�].������}!�I�֊O��ɿ#.�Mmz�˭�M�`�<.29j�+��3�i��
��1t�\��]{w�;��:O\�B�^�*�Q�>*-g1��z����5��L��8Nj��%l��^�����΃����xw�zznWy�03V6��L	������V���\y�оcވ�b���Yt��]̧�r���I� ��^���L��E=V�#QFiT
KP�%���[��?Gjys:4%-�Y�N�@��&� ٿ��d���#=^�
�qT��Si�s�Ǧ�o�z�h�����[��S�F�ky<�L4���{�=�>��%17��) �P�Lco����hc?��?C-�mpߚ����2��؜J`x�����#2��.[����
բ+i��.7 �������Qs�r��;Iě��J�����[0�k�u�ų��a���g���Y��N����%�vs�]Y�=D�ʸ�H?���w�5�7���|�}.�ٲ��y���ӽ~�;rd��'�Ƙ+|��k�\��\��!?S��^�MD[��)!=f�D���r��^�'�K��,�]Ч�ۦ�bU���^#<�3�sy[���
�n�҆�,k���r�ɩi:�=�֪x�&�Z' �7��p���QO��v������K���u����ȴ���p�`�C�����]To�ԏ�/q��£7h}������K]-������*RH�B2�|+���ŧwkw:H7�6�d���[9ٸ�� �����R��h�j��]�$U�8}�ɏ��ƌS(Gc�\�ͧ1kU��LjWI��YJ�A�[�އS:��2�-�~�0�����ܫ0����5�Kq�����E��>ן����lT� )k�7b;O�W���Cz*&�^����u�P�$����Nc�}a����F-���=��b`�$�m��q�U��:��|�z�ݵH��P�#�F3+�Xjqb"M|k	�J�7�"��Mq[}K!j�U0��d��g�㗰�K��UB��,�,mCt�jy�~F1�n�Yg���Y]��P뒇���3�ΣC�j�Ԭ�Iޱ��Q�qSb�������ц.:i��bu�}�[3�G��Lw��xۅN94�fދI#ʅ\d�ۚ���y���b��.2.��	M٘L%�p22�W��!0������@ޝ�j�;�ʡ��8�JC {|�c�k_����9Β�����ޭ�_MB6醛���s]��6�A��%/�)��Q�/iZ�'Y�e���T)e��Y�� ��-�l>���!�Vt�V�s�?�l^��!g�os����/;)�=z.
���N��o%dA���<)X�)k�b:��<FP=H��ؐ�E�g�d٫�|C�J��p����F� �'�����|}�UV3oHRU����B3���'֎�-��?>s�%����Yk�,�E��{/�߻�2<ɳf#�����b
�k~x����4u�B��C��ӌ|�-"�?
 ;��]����������V��~�jB�#u����ލ�b�Z| �� �m%���@U�4&���������.7��i���@����ׁ�P�ff����(0�Q�_�����l�Ҏz>С��n���%�[z!��I+� ��(���84i����"�Aݩ�=R�*��1>�i��Rg-{�:�H�څ��e����z�d	�-�1��j	r��j�x�8�z'4�B���d�_C� G�{ki&�u���M�𢷻���;~�������^�v�� �+�û��럇��0(9Jv��h��f/r��Nr���1����:8����8(��K���(�y���ƺ�x���`��0���wvH�/���gTS��85<�N��ث��7?��7}u;�{!伖}�z�!�x�����ֹ�1r-ө�� 8*��R�K&	q��Q�ɝ#�'C)����q��<1�	~eݠ3|%�35��0I�8b���U����eocQ����h%%���f�0���3��t��N ؘ� S��q�ңT�݄lS�Z�}<O#����w�?�3��a��U�;�r�r��.�%�1��4�h��Э�!�p�o��=�7	_R�UQ�z�:��IlL�'�����h��4!�-����u�L�1u�ߥw/���C�x7&�@k�h]�jYY4 ~>L�yS�|#l{C���V��pJފd�q�Lʻ��$OX�;u���ݩ�#?�3��l��7�h��@�\�K�}��yt���ܲ�!�]wm�;M�>c�B>��п1o"$&<�U�2Y�����y�I�KT�xg��j�u� �B�^�Ww[	���m1H��߹AN����M�.�'��%8K�����s��<ʴ�#�<�*/����U��h;ȟ�h�a��h(8Wd�WH�&�����tF�v�6�ЙBs1��0W�6܌T����}�
LPA���䉺�A������`z}Q���p��-�
�����b�|a����{��;��F��wF��je	q�.=�G�Ȏ)�2��5�]��p�ס  Ms �3}}�FG��j�)3���(��w�],�}��5�ƕ�ݜ���J�L}��V����GȞ� �ty�������� ڥ�3�"?�B�V��7���]��6y
I�啄
kPɸ����=�x�:������s �~���x�;�[c����_���W&�w+&��\bۧ0�h�Ή��n�˝����̛�w1AJC�y�!��f�j�&Q����P"elp��?��i�2�F��f`P��S���O
cZ,W��_�8�8�쬒��IÌY�{&J�	��4
w[
=sXzIk���c��Wrd����g"���D4ɽ� )��wxa	k��#N�"-f�8����@�bj��K�X�0M���a��-:"�O����B����ʝҍ��p�Q~wr���X�%��K�`��5�^b:��G&�W����S\���4Xka���*��`=�7ɰӗz�^,t�>I��;E��X׷F���uN�0�F�@!�v�`���j�&����,���<�M>3��,>Gd�x�(�u�'�R(�р�f�SU*�kz(�b�4���C�}l�$��T?��\�ZKb���ؕ@�C��0]�7	�t�f��9�����?r����K��V���a�o@7㣻Wc*��E1���v�м�	�s4�\n�@�=}���/�]A ��$%����B'��[���QWy5h�j���@�H�)y�!��7i|�:ޖ�7�Z���N��"�m����_�s��Q�{B;��l�2�(��S��i����4�{^ǅ`�N$�Ap�VB�X�����#ɮL�>F�)�r�.�4��Q7�f��x���F\�F�s�l�:�U]��ov�	Ӎ3�N?����߹#CQ1�$`/pc�^��;���G���T	�
T��&���,wr1ø,��7_2H�~�z��k�fF�
*~Ģ���fr��ъ(�z�zO���``�}���s0�m�d&��n7�K2P����~8��D�@��/��`� �� ���H���c����PB�j��YfX�#v���X�V�Zk�(��:����C��f ����4v8İ�t�s���OEw�[�����Qb���_�jמ��ڤ?hr�Na�r�����;�*]�mNOK��O�n����ܩ�YC�,�3������PU���a�D��ѡ��oU�$��ΝzZ�Z�^K9td����4���g2S�wu���^��}È�K�%Pg��q�q�@<��y�F���=`��N"%Kr,�=�,i%"�p�Uc�4������	51����G��@L�������,�꜌�TF���Ӗ?�ۘj��Mp���T<�,���8���Qd��nw�~Uvu����2���h�߱�x��0�8.:bK>��Ć��[K"w�8%���u3��9�+6�Se��蹩d���s���*��������sI�C�j��"Ǽ?3�W`?gd����U��nw���%��>�H�����z����� Xa�y@]���˺��-�>y��ʭ�>.nQ���l�����i�pl��Ԝ J[�ho���9�	�d`yU�x��Ća��+�d���-��>��B�EM�����%@�Ą�@���(�N��E�|'Y�5��9�D�:䮌n�=q�8$�4��T��Y�eɱ�b�O�@m�+����|l��Z6�c��`q'/栴�u�lr}!�#���Z���y�Y�V�r��s� M5�k$'B����C���L�I����TNH���z�Y�Fβ&��uhR�����u&��N�M��q��+���1.�K6��57�PWs%JR-��3p%�T�Mg����&���ޠ-�?�Uk�E��~�b�֗����akZ"����vxN
N�����Ls<H3����+��4~�G�߁%Q�g���^}�fш�z<�͠3̱��B�-5tl۳<�zj�r0� I�X1�yJ9i�<�w��5^��$!P�p�A�Y�����z����Jb"\3YH�Ǌ+��
�Gf�U��;y���NQ�~�3���"�஽U��K+S��?�P�5�j@-7T��]p�"?�d6�-bk�V'�,9�����hQN��\K�oF ��@�$��\�,Mc��}hkV+Z�����.��4�s/�����y~�ϟ���X��6V>�.�D��> �_�CؓM]�$�Fb���w����݈qk.Z�H�T��]_GM��g�����E�|��^ի{�(HfK�6OT�M0��wR��K�]��*\�Y�w�G�7�і�4�ο�fIcΞ�&.�v�fOn|�����O[*�mX�b�,N�%Ƣ�H�$�d���\���%���� 4��B.�y���?�9�������0�)���M�9�u�{���`��QkX�7k�_k���G��Y!O�oB+H���$��YV�]��S���A*Z�ɗ"1)2=M���_�X�/�xH\�  �;�i��$$�w�Y֞���*�}�̩�g�t�<%\��莖�U��@�&W�'����u[�$;�"�ׁ��!����)�	��R,�n�[��z������z��
/� �����ZK�~:''%���=2�/gƦ�^IYd��[����eL�A΢�O"�	�c���ȟ7���a��i{ǯ���l����a+��R�c�ij��Oĕ(���;|���JV-ߛ��:�ۗ��աV�^�cv��pF%;M�P��,����5���A6�h��h���Ģ� ���U��4p͎�%n\��k��ۋ�^8�U���A>�/�����h��k�0�5������a�W	M��T%E�Em�a9��42{ ��9����yҚ���!�B1��,kt4�]�%І���7���1�l@-����-c=��P����}���V���$������ɄYL��k� AXY�g�X?�P\L�8�	�[A���4W��9y/l�j���uc� .��D�y����8��d�ޝ$��ZTe8��&���HG%^����<ΐ},�G��Da[d�@lV׍��a��A�/��IdA�c1�y�C8��+��&�r���3�!�#S6��qB�G���n�|nG@6z�YГRm�l!���;N��b=�FqT�r�Yd�vA3
�Vu��.sJ�<�hi`���_s��.�WR4�`h����g����8J��@8r;GF^�;S���M��|(-�䂱u����8�K�B}M�S���T?.M��ٮ��w��S]�l��KTu|D'^�9nm>�W�����o�TF �������C��lP]�4���%oV�+���ǈ6F���{���r�B"3���@'��{�<sjT�4��r���1h&�Z̦�H1�8[�ʢ�[P� h�f���QX��,Nh�֓��[��Ci��Ǽ&�NI���-L��V���h���A�U�˝Mdy���
�Z�~���y�gV=5��`��l�;m����B:��e��e���@"��U5
Q����Jz�󼬫	�s&B�Y��*<��O��@h� ��nzk-�����L(Lj�x�N7$$��F��]')�_��Bʍ��P�9�G?2+�1�� ����&�)V�(<�lP�)�C�[��7��^���1��5n�FH6�'��G��:�}u�8�`>��$��q��5�zj�s��%��>�!�����:��8�S�L�$��2�70E�'��3�"�̪�������hZ=>��\nf"���_�cN���U�D���@�s�
ƣ�]�!���"v�o(|�6R�t��D���v��1���<��ul� �����ؤV꣉?������I�Y!��-DaU/��r�@&E:�u<��6�R)��o�4��Ӷ���h����f���9��,��Ձ��L�G-˯m�KӕɈϾs��f����B�3m9�;<���R"�˽;s��e(�* �>0�G����mrn���g����VBO_�B`���h�?#
;h\�i�j���=|�7����y�b\}�a��# v���RT��Dd5�.F��9�ow�9��G�h��'x�r�����Wm}�l��6?1��<6?G*{��V����B�)��h��ґ�^z�lYsb����W���c��Ó���T*̈́�Ρd�t����P��U3���rS-fv��X���!g�%9�����dP����vk!T��k`M�J`��E��q=���.����M�չ~h��T�d�Ki4��i�,�4�3�74S%��H��dŶN�(�>w��M��8�K��i�n��3����}yU��C[����(
�O���H�	Qj�%KM\ʚ�!}��1���v�!��ݭT��?��M怪&3�+�iI��`Ǌq?#m��mN��g'J�W�u3�=�tGҡ�Ѱ��%�i�����m�6���L�'3�d4�ѕ\�$�`�0�T�O1'�\w�N�:�b��7�����~���:Ĉ��w���Vd�)�p�k$].$�w�ҍwR
�=&W 2�1{m��Ipn ��	��Y�&t.��Es��C�%�2N�ePzQ[4�6u��O�`����<:"u�g�-i4Q~�˖\P1\U������N-� K�+��V�u�4�؈AW�b�"�v�3��$A,�4~�Ch�����Y�Ĺd���P�W*w$|��	2F�"z^·S��]	��bg������W���9�ڕ�H�����_�2�&�$<,݊�b9욿)O�	�_��^�=��k��M�O6��Z!6���uN��y߳f&h~ ��{(���D�F7]�s~lG.P�́�cv�v�����i��8��G�H#$�7��Y�_�7LX��-��8a�����O���/�����hJ\́�$�LBO}N��h����L�1���ֻ�/h��]��Rn�nN�7p��l��/��p����I8�8�11�X���\Zj�C��Ȏy7n`��ϖ
<�O��t�����.�8y9%����iP��Nd�Gy�B����~�~�.�P�(��.�\�sc�|g��_������ k�P�3L nQ/��o�v��C�c��q�g֪��N��1�f~��j��꠩!��<	�
P:d2�C��A(�(�n���x�r��^�+�-y�_-�͋�2�m" VI����.�|c��K�{��Z�MB���X��q۪��ؕ���F
��#q��C�7e�a��݃�T��J�3A��B��/�~�$��95��+�墼����y ���B[LD��l��DH�۬�f�V�����LH2� �LM =�����r������x��1�MJ��9s=qtƇ~!��=.�7X���O�-�K)�(P���AƯ�R���\s˭��֖�%����F�Y�*/"d�P��0�:�ȷ�h�����@���[�+��?`l0�p	� �mќ;��ō'���MG��%D�:AUL&x�vM>A�; ���2�$�Xҁާ	T����D���\�2?p��(C�$2n�&rY�V��r�gTk���̧a:�-*
E1c��F,����+2��ڮ6{�x��j6��71B$ +���7��uo�l �Bi{A���O�>h�C��jg�/Q�y�t�s	��UZ�
 ͺ}h*����㥔 �pr��>�{<��<�c��ۄ
�M)�H v��&��u��v{S}�|K/�CiԫbO7�#+��O�$��a����˩�j� ��c�]6�v���l����'��'��d!����������5��2��X���Sr�$�ʃ��mV�2c�k��X9�;����X��n�:gt����+w� ��k�K�5�l��A����#�F,��Ly�:W�%��Fl'�k�F&�N�k�+F�? qfG�h^��x�B6���%m-���/�V�1�eA�>����U�:���4����V�f��n�_&����3�/M.@ëq���.͔Z/w#
�P+/��u�����1L2��t�׫%�F��F,5&rd� Xkc���V�!'���/@1���gB�Pv�a%�\[�6Q�z��OFG��f�c�~�W]T�	f@�fX㔖����pOg=� Y}���Q��WM����R���ہ�x��P��i� ��ۓ�����Dbu��E� 3Z�A8����k�+��h��}s��r����Ys>�!�`q+!��Y4�D�q��8�U��e�����W�]��$�9f��i
j�@H�$�j�x'��Wm��.\�����:]oY��K�jD���ӝ5�sp��Q��wEu%��ʚ��'��+y��g�Y'�b��hٸT����Z���촺J&ſ�2�WO4D�eX�R�Q��!n|�9�x�A�[�;L�@G#�lʊ�v�w���s f+F�ޢ���_O)��v��"��Fa���w��KXں��L<]*���{M�'�{۝�Nx�狼��ĮY3N:�
ߕ��p%Ǟ����[���cx��7��t��g],5��{� _��r��t{,�~�V�R�G����ӧ5ư�sI#�9��RȂ2�hG
N���*���B1�z1�Hх���)����86�1u��^�y���4���q#�N��}6��d%�����{��X���`���|3�V��n#����<��i�#�[ e%\N�.�<�KL����`�M%�y�1n�i�����B����Sd����1Vy�}rS�9�&��hb�r*���R�X���
(�F�I7�
˛_�O�U�T�MA䷁��N�;��2��pU��H�\�� d�Os��QP>���rzw��JI�vA��rqN�ί�)���D��̠�mǴ�^��w��3cX;���WjLh�8☈�x{��Kc2�Ǝ+�ɮX�ɤ�D�oY|��TI�N���>4rVx-�{GH�**���c�3IAj�um̆^,���?�$��ϡӥ:�a�����E[9�A�n���%M���l=�b���� &F�On�e�xN������(��۫2����/riy$C�ν40.,_fn�؊��b����&�<A����#C��A��&�h�޸��p���B-��de��db'���\�q�X�gyнm��Zy�u'�5��⽇[s�ڨ�����χ�y��VN��ݎ�
���p���U;L����Ve�c�Ɍޠ$�qAݔ➎���X�5݀MCi��$ϳ����T*x0�s���k:o��������̧�|��O��A��֊!��ChQ����3�a�*���b�em1Wi��Q��O��U�\B�FʙRl�Z�8��mp��傞�"qv�m��X�!��0��D��Z�s8���|�a���6�eR.�(�xP��FF��=�adl�l��"�t6[���� 7� KL��j�kv�,M҂<��
vG���,�Oc`ZA���7���d�#��-1�K�2�sM&u��*I]֬�U�%K��#�����ܑ�<3��zd�����<�xv5b ���>�TҦ��9|M�{���΂�rr���P�s������Wl�l,��Kߊ�R����[�鉑��@0Ȋ!�,Nk��R�'�����O)(_g����Q�WwB�]�wqʰU�R��e��i��7
�'۳��C<��
&5����4�r�o�z�k���R�³�����6�#4�aj�xAe\5a5��߱��[���i�Ȣ��;����x�@#�Pa��V�JJ�K�G:�!�-+�zx�Ƕc|���v��ɛO�p�y5<r@n�1��r+�u���QdF�C8wS�h��%�����55���<J�7�S�Y�C+�)����h	���7k{+��.G��������R��!���4z�C�=�JY��kVЃ��_4� � �tZ��j	U�/�rU�C�W��E��fK �5v��1+�{��V>����j�Ox�%֦�6IR%��4=5i��t~�,��ލ��CȪe��G1�5:w%�F'B�Ú����w ��''��rJ�$�F�Z��(�K�!Wh0z�CV��-i�����t/���,��p����vB��H�bV�F�n���d2�����ȅQK�TPz?�x��s�n�>&m��F���)W�����a�vbrDI@��*��P�3&�O��nL���$܆ �Ϡ���ͼ��jK���:!HA��%{�yK�9�����^vnty�6�K?�dB�I�	}{�]�� ��p`���E+p���V��960�;�G̒��i9�)*��>_��2�a��?dD
��ҌT1%����b&�ď'}��MkxK��Ql�Ԓ�ڀ�x
�- �Ǯ�o��Z���QM=��0fG+��|�k]j�o���sTC�4:,Qs��x5[R�ǻ w9�4�R ���lD��Uf��[�!g�"%cb@^�+�c~-Km���(l�$J��!�(d(u
t��ՍU��ƣ-k��}J�7D���V�Rҭ�*��	��ˏ�I��"�x^�1���$Xs��u� /�z���ٹ�.I� �7
�r��iiS@�ߏJ�F򛋬�}�f4����y���T/+��+����_Qz�,�r&9��Q� @��o������[m8
�yy��D��D�%�#l9�|�)��$���RМ�j�+����۱�P1�8b_�W={AR��)��$�Ce�9�?��oC�sT��zm��Ћ� )mVX*��w��nqa~J�	f�����Q� )����q��%����׊�����:%ʰ��sml���`~�}���o�&I����Rx$@�/2i��#�9z�>V���ڇa�� �kX��ު��+���\�o�C@#�jXl�
�.�w���v�K'|v:�$�r�K;m����J-�l/����S�Xbl�
��s�.õ]Ԕ���d0n����*��MIg�j(O�c�9ArCV�=OJ�ư2䲅�L��|�70KMB�����)+�(*ܿ���@	��WY�w��(f����XN,�S�>����n}����6_@$���)�QС�(�Bzoq�MeA��t���F�*����ir�.'�e��>vh9ۃ��Za�����r��FX����������/�����(]F�	�ſ$���w����c2V��n�d�,]�wD�lf�L�W��(�I�єk^!.���_\q5b�]���<�������l�\��+��eҢ���#�n�{��;~�������,t�ǌ1�ܕ���P^;��r���W
=3�ZR�bmy��m^�[��>��� ��/�P��ͬ4%��a���N�!jY�6Q�Q��b������L��6��v����G�6��W�R�b^��RMžw@ �䥡0�t-Gg�o��9q��t��-�%ߦ�[��v	؃V��=�.
D؛7���z�Ŀ�I��n �J�� �2��7B9��~C���VO����xɌl*���d���Mp�g�+2ޅNvou��.?��R0P����H��W0�m������l��\R��.�X5>!�W�}��i:���Ѵ`-1�=�^}�/p�6U�zp?z�0����UE���b;<���h]}B/妩y� {[�{�&��9�/�D֋�	��"�H��\|N(�$Mϩ� ����W��?S�_�k������|�]�T[��7mv ��)!�^�i3#�|G������6K��J*P���s-`>�Иب�=\�2 ����:��!-�Bc�&B����p��%4-�n�B����B�N���mi5����)��sc��B�09kZ�W1t�D�|�����h�'��RW�;3��[a�]%���쉛s����87���8XRŏC�'��BgA:�wy��a���>x[ЖO�/���u�ߏ�0i��:��1#��-�;ss���+��=����S��´��/|�%6	��K'��Ħk��8�(Y�,�%�T��l}PN��@��4=|j��Yk��a󑼬����f��!i8��OQ0��oXp�E���� �$ `O�J
l�W�"����IO��Y�?R�)��-E�� �8`��F��niU'=�"�K�pjtEˉ�k-�-R�4��3C����{�0�g�X	bL��e4���7���:B���O��~��kګ����l�*�.����7��q'��J�RZ{m3+�Ɣ�^���*�r��L��d~э �c��J�e;��	>j�c�����F?D �	 ��ȍ�jwWʾ%�_~WkC�?���}�Nuo�)�5��ӝk��'U����8M
��Lǩ>V���^��
d\�KX7�t�C�� �=��s�&'�,��Q:�!O��둖���d��W��rt��VӿD8Sg�7瘟QHؚ��Gb����1��r0�F�v�F�����j'���M-������x;�M�48zK�M3����c�N
���U'�V����E�Fk����+]5l�� �ON�I8��)\��GI�1�lx�V��="����������~�)b��{ZE����m��/�7�7ͧ�>h�ƌ��O����)�y��l�oX����>��]27�@L�����h��06��*B�'Pb��r����!��T�Ƒe.�<jզ��)���g�8FxK�5\o`i
�og��,�`{VQiXF@�Y28ʜ�ڡ?Y�'��93����P���;X�j�U��D�#��MxZ#y��.COo�8.лk�I�Va�\��bg�6�����9�=Zj[�r���7ݖ�c�j��I=���9�?�r�;3H��v~{� �A� wγ�8�V��|-�m���L���	�Jb����%�{OQ ��^ޱ���t3`+�ɣR n0�7&sj���IE�����3!� 
\�h�^�[�	k����0�޽����Ѝ�/�� ܤ����Kh�K��hN�>���9��2�+�F@0�L^Wƪ�$G��H�I�o� {k��E��(�J
��#��H��i�[�9~'D5;DBkja��s/f�a�xń����ns�p0�y�q��C���6�>B
'%<ޟS}�o�Y2?�\�f�c�5N�����94\4d�t��g�-X��.܇�;�f�O�7�\W)y`ȸ�'���v�L�Y��goN�W�����{�$��
C�����jg�H�$�/�;i�a���%���.,��P�ctG�{1�5�`��%���wפuOf����c�!D�9�f��Uc�_NS
n/9��>�mѳ�+�~��0Gz�1ٗ���}w�t�4���i5�+�YȮ�tx��JO!?�-��S�*(���*��p	�8�)�=�+9�E�����Y=����Cِ8ѐ�Gއ��N�8�5��5��Ck|G����PӺV�'� 1O'\Jq�$����V%�a���F�NK4��Ӑ�+Ia$�0Wm��Z�s9�������a����Aڲ�G�Y�H�f��ⰵ<O	�O��Zգ/�����Xͭ�P�C�����r<VI��ޒ�A!(�]�$����͒^�@j���6��+f�0|�nZ�'�H�
V�Ƿ���S���n�Y�L5�T�����hG^fX�%�x�G�������qN��#�|��5��Q�Ǡ9�V��
�q򵖑Їuk4�"��	X�qW�l'����κ�^�M:v���C��zB�٣��a*_�[���@:(�.5!��t�o;8���.�Z�=�</36EF��+��X�Mt+I�F*�x�^0G3X-6�c2�X�Il\3DH���s��K���D�s&٥h��X/Kɡ@��o�H^�	�z�,��G�W�@�9~h���(i��n�m�b�e��CI��%�5�$�xУ԰�k�F��S��A�a��J�r��ƌ��0x�˥7ц�l8r��)��P�,�;桉�l��xF6��롽�Z7�	"��Fٻ����<MG#�}2�H�h�y��k�>C��4+ާ�Rc3����P4��FHY�,X����ϱUK����=fBYaȦc�6������m݆��|����1�GT|+�{3�q�%N� ��*ڰ� �N�����(�v�i���v�v�#^_�!�?z.n�-:��O��?�6SKw�k�-���Y�@	�ez����9IG�"����P��wӛW��@��2�a����~�f���+�G�~�?
��Kbp񭞿��h��2x��:m܆J�>3o-�	�Y�[���`�1K�9 �,��qx���#`9����1�0p"!��`�/v��O�%�J�'Z�*�7T����G� ��4j4�� [䤭m��j��x2I�?�W/��V�"�cw0�� ��Yw�'���u�B�+�n�J�f���ȃ�.�ב�2��÷���L܋P��?�^�&|�'�{��wz!�1n�\iL�cpcu�
~<7�����C�m.�9n1�6y��Nn�>�c�g��ҿs/>[]QW�Xt�ә<� R��h�v�Q�Ul�f*�;�h��m�����(ş�K��>�1�h��V�ʃy��bu��s�'��%��N���d"Wj]���
dǆ�%uug�m�����~�u�(��Y���i�s��M��u*�72g��v�����?+����K��/HU_�� �)N��y&E`�L�*�=�T��J-���_�iX DiaEs������fr
pJπ��#Ҭ��20S���e��"ݐ���� ��%�#��4T*T��"��j��Us'ǘt��B�a�D��%�p�'-��9n�|�ۨ�U����tY�z"�˭]uS�N�of!�S��m�j����[WW�$�KH崄�I��ڄ�`���KD�׽|��mM��+V�d��vi�6"5�\RFx�=��������jF�}+��X�5!:�YJ�ӧG�s���UG�����.8w�c0����a���ɧ�Ro�n����ּ���1�k_)�)���~r�j��~x�^n*�o~ڌ���Q�\�w�|Ѡ��If[z�P�2���
(���bǦ��u�G28a�3E��_�/�ȸ�hG�&�:��I��Q������E��^S/}�S�?����0Il�M:\~�'��M�#�I�ar�z��O�6�3gL鎬?��Cl�P=?�f%`��=�[��C��9�9{>���L�^1�͹���R�Xt�K��'5��P�8��B"��5c�n�^yz�q�U�v�̒��(���<X��<����:���#ه�J���c� ��zc�^�_��:r=���/b���f1!�K�vB����T�V)���G�̀�c��B�n����A��RD���i:�$�X������,�V�~��]4�"?������m�J��@�lXk�j �v�b7C����Y�J�ߒ�*�O)%�^#Tm��P�Ϋ�3��V�WcH��E��b�h��9	i;����)<�:�'�"}�v���
2��#`uQ����� �x)�m	T���<�h� �"S�4��c���3.�����4�<�����D����z7��C�7 ���Ѩ�~���g�g�: ����p�D^�I(�Q�&g���g��q \a�75a���r���(���骁�ai�2a��-��5u` �ߎ;8�n�%#hw�c,��N��ǩ�4��%���|��Z�& R���dπ��@����o������k����iBj��LW�ݶ��E����GZ� @��V㝲�=O�+�x�hcT��7����Fk?Z����}^��pҕ����J�p�L%����lzD7���,x��t�Ƞ�� �`'�A�2J�}';oy�Q����*�����:����F���8�3��+�<z���	D���������z��$���-8���N!�A�}o��˽"��p�v�y�Z�q��=����3#7G������o��cU�hX��]���2��h�C�a�9f�yd�F�P=s��bȓIW}YG���_/�o�#���	�������$�B%?�ثjo��6���ܫ/$�=��R���`_�a��1�x�j������&�]Zi��4:o1}��f� B)�NEЧh�՟�B`3�9ؑOT0Ҵ"@Z����G���Ddxp�-� T5�}�g\sB�^��.c+�SP�VS����!�/�ԈE���}�qW�X�"n~M�$��2�@���H��]C�$OR[��֑�9���T�2�Su��?kK2�jDk'_):q�"�w �4$B�&_XPL��j˱G�����oQ�/�EP��xXP��X���Y'3gYJZ6�,@	�.�-�rH��%{w�>�'��ՊZZBg��t�@k�
���I�\=G��bQf5UR�U�Y�D�@�1�?����l/zoI�ܬ� �q�
p�~%E'��M�GY<��:,A%�}y}[[����$��5R-J�m��9,Ӄ�yۆ0��U�
�։*%�x��5����z��~�ܡ)0��^�S�Ee�go�#p\�cKm� 9�Sk�F���{,G�.5���:x����E�@�h�v�������7�$�j�o�q��};A�R/�����K\f�P":��F /T��Ժۧ�!r�9n��u��L� 
Yw�lp�q ;V�a9��
8� �N�!f����.�����k0ցM���;O����i ~�w����0���I-�T�,i���d���4w�Dh��@��,?��G�L��{��Ix۾����撴��l�Y]��
�v�9,�[7.��tw�n��W�'�� ���mvW��y3��D��~A��Ǡ]��A�h�N����խ�: ��l"ѳ-�	�*S��$�y� �͞ԡ8%d�:Do� �s�`1�b%��v ��z)+g��k�iT��^yf+�^��Ʀ:��51t�#]�5���6)�`��F����J<g�7��������*i�Y�#��Cq9���Z�DEn1��yI}.�0���1N�eG�YZ�iH�g�_Ԧ�� �#��1�&b�O[l��9�d����!Ξ���>�i}����^u�����>�B$`}��T��t�>�9d��_���O�3<@*�o\h�E�'ǁ��B
%=[QjZ��vz*P�*ǡ� =\�R2�Z�
v7���YqH��PY!\YW5��&�c�<�_�نp��Hǣw<h���T�$��@�'h.L���mw�}����e�!�{���]B�Cs�q���nB�\;��$�A{0��,[����4�	>N||���v*��L�����17<C���i�S����g�<��,^-�)�����)�V�λ��CA��m�M�R�(�*�l���0�X����F�q��}������MNӷ�Z�3tT����(�}* 9���t�Z�Ue"����.Q�cS6[M������R��7��PF�/�%�R�����?��(-��X����
ZT2C)6�~&_�c/���1 �{��"v��9=cJɨ6rg�6'm��t�M�t�}}I��W���V� ���ͫ(�먈�T���3�F&/��#�Sp�>6>�<�ec��D��ܶ�Us���h�D)���mמ8�nt�ݟ��W�hfux�]3G��q�t��#�b��&	e�������+�OL��}�@�Z���J�����:\ߝ��Y-2�8�Sfu�vħ@����K�l-U\�j������?���D�]*Z�h���`�B�����)V؂�����[���}�BX���+�?k�SN �m�/(#���IR?�����t~E♯H^���U��O��:�~��pB%̯����:����K���$8i�m�!d��<�0f���_w�tX����]���<��:��eDX��н@5�b0!��+z��iƜ�α����~�`�+���Q�)ǥ����!3r}aҺ�z�aĞ"ү�n��Y�h6_���^H��_S{f����a���p�y�A��3�^�[�l���~���o<�z�;�����>�g؎��+ʹ��^���_��@,�r>⠖�̔�篜/s,`˵\��+�(�eO|���4z
HϺ�kڕ&i����ӓ�.z�νN��:��2�l��+�"
�R{�ɝݢ��~�6�<��ʺg����t8.�fhڑ:]�¢%-��_����7N��i��S$�q��.P
��.��~Gc>��D����߿��Ƅ<� �zݞ���k��Kzm����:��=��tj�b���\��h�]LMn�K��unn%l�;*�FV�đ�ݒ��.��j��x�Z����Pw)���`�2�5��W)K�I�! o� ����ᷪ��]u%@G�2Ď3���bތ	�h��:X5��	����仭]	��)z������,X��tJe�:���5�&�y,-�D2��l�x�az��7=�TZ�mR)�EА��QO��b6�I�o����]�r�QU�P�UX�	����/ȇ ��c��{�����ĝ�908�76xյ���m�?����r&	|�jNrCx���򃼔�__���z��+�%�K�����z?6��	MסP�0���{�1�����Z�9� @rơ霊�F�Q��+{C�끽5����z�A�w��)`��4fP]�A6 =��n�24Z?�E���P�t43}�R�{�~P�:�D4u�$�9�$�={'��5�0?�L��̢����艓��qb{[�$��8�;��/
QB�7Ľ��g����GF�^�,� C�[�|m�U�\�s�)��B>^��f_{=ڵj3��l��Aw�dwj#.�G�ϽB�aYĭG����2�h\z���獢w�
j�(d��y�R(T�	_}>6[�4Ъ�����?�|�Z��'.�Es��tۜ�$#�k�ӻ �+�
�_yj��T`?ӝg�Mv�Z��'F�|2L�$k�>�=o@6Z�x�:����+\T3`:A9������Z��6_IJ%���}�sJQ�ܼ�A�r�����/�:�L�d��4��I�ex%^,��Ѻ��-��.��_���n�wi�v��8��΄�����No�_�'����g+�L���IBZ������ϸ�Q���ہş���P7�Dd䬪(꣗��)��{��Ļ�Ԅ���H�l�ʋ����s�F��A�xzl�S�V5�y��]\b���S
���M�m��l%��=�}&�`k©:�}\̜�6�w�ҎBg
��F-*���?���1�C�W^�E��o.�뮁��D���L��t".�D�ަ���KmP'��9.l�ׇ�D	J��>U��g(d�u*T�jQݐ���ng�������ػ�rcQ�3��1�gG�T���\�f�a	�(�?:�84VRU�ԐH�W���6��ʲ?���e��,�C���J��ǜM�m>s_e�W���@$���m��z}�(�&����U��z�w.!���γ�d�[�f��s�Y=�!m��[�H��^�3?�-c��K$��B����kZ}b�j�a�f���꣖�(c;E��Gw�������3�I���Nƿ��[��9:�j$K�]��!�o��7��c�q�P>�s���H�:m/�2�_��F�l*�h)ǰ;0"��Lmyn����R���g�����d�S�V�+���|0�H��\�5���qGr6s� k١�!���]�_M�n���F�2���䔀���~9ô���h���e�8�o�u��k6B\3�HEV7�͆v$�c�x�%���4�+8�����w���	�/�G3�<V,Y�͐k��k�օ>����܎��K�j�<��*<�Pb�Ǌx(*!�P����D�$����}+�֏���(*�m����*�g�
Zw N]�
�ʚ��>=Z����Y�#��D����HC���Np���r-OO7p���<�J�HU�#��k�f���p�M��8US� �.2s֫E�n2�M�Tٟr�MK��P�����W���.����d=o�v�𸔉�w���Z2��c{[����[5�I�)j(��)�]2���x�u�boB�eY�L�pI�{k	u9Y������{U3�"�_3/���MC��
�n�;).z�����sU�bCZ7�Q"W��C%���g�,|��T���i;M��I�IX9�Z� P���(ꑧ-�D�J��U����H'Ŕ1)����!<x��G��;���=K��!�������*nm�f��%eA|ɉ����޿4���A���%4ogs������ s���S(*��wbw튬q��\,�W�
�ƈC=U�a�ե���d�wIA_%2O��� Q�C�w[�|�V����sp������"�����u9�[��%˯9�vY�a��W�JP��b$+'w?z�2n�^}c<�E�f4�fZ��B�z���vO�O,|�����"�z�Y5�(�n��	}M|���5�r� "�z�2=��B�*FIq�|v��6�o��i�H��I�-��Z��%�c���|eV��r���\+���n�aI��{Eo+��7��	-�D�2��(S˨ԁ(�	��}��i�&��s��C5����`��,�DB�v������{zHkU�𽫜M�,���:ޗ܌����C�t���� W����۾�m��   vud�x"��A��>,Z�1���j���{#2�'���hd�({y?g4]eȸ#(�9�m]��tZb�+�.�#����y��eg��k�Z �;�����"o�'/+j�gl9'���/�&��	�8�+�Ѝ��U����+��<�lz����a�cˏ�!�Ł��Gx6��G��)�yW�e�ώ<1ao���M�p����[L�^{����z�F	��`�o���YS��ji�p��9�u�;���y�`.���|A���>�َ	ER�b�P��6r�� P�H�<)�|��Z7�����N��I�ї�-Њx���ͭ�װ�ZQ�F����ǧM}n*l��y�,�!E4|ov��>�~�zv�wS��`H����$R��iڼ�["�k��F���M�gAݶ�뽮iTӧ�x��	%�J���&t�>������P?��,��9��r�k����waq�$�j����3рҜ�x�ʀ����Z/�˱��8�X�Ϯ�7��0{�֯�8��Rs���5�n�F�v�������7����3ڙSP1��H0�d��F�I�7š(H�z�3p�e�M*�0b���q(�; ����]�g!��m�N_TJ�kY��u�"n��x��.�o�w��eS�$T�3�����+��/��:����良L��W��`?p���\���Z��`��p���]�# �ŽK�F�uh����&��+��XX�����a�U�U�N�1ɋ[��\~�҉ǜ�g�Y��S�e�@H
i��3w]�t\.��I+5f&�&(�qJ@d�$���R��4��'T�	���fD������4��MKVX�O��䛕zj��-�1+Y[ �2Y�R5��M|2"+o1:��P��xe�A�'A�T��Oゲߔ/
���������z�
�A�r���<=w�F��p"�EBP߂٦K�:2�T��4���`	@^yRJF��]�p�
摯t+c��kCG��:�I�\˻��h�#AY���q�Z&��J-NW��49��,�4�������M�i:#��44z���!��嗡7��p$e&�.|=���P�b���ѦI�]�p{�q�X��"}�6�b����[����(����Rv����"���o����m�N� Y��s��[Ѣ�j�F��u��v�G�^���ty#0���}i���� 詸2��Ñ����-=5 .Nk�b��Sw��׻۩H�Qld{�4�di�g�i"�����܍�r�\�&
��Q w�.���.v�g&�Fs%3��ź�C��xʖs�x�Όd������`�?5��p/����*q�8��C۰$���P�W����e�C��/�<�ƩU�7z	���c �v=�C�L��<� ��($  BEg�ǈ)�|1XW��KT��a&x�!>F[gU��O_&-�^�Q�w-��X�!lD���$�ߴ��gmGy�:����8:���' �4��Q\q_�*��c��6�s`Ǚ�bb��dֹs�Z@��W+���:�M�T����^�q�<����F�Ee`���D�=>-os��j®?(����<��\a`L
=|{y�r`���й5E)�﫱'���.9R���g�8C����O���qk�5��6<6�� K[_K,e�g��{���S���n�m"�ޝ�'y����?�h�^�;L�>i��29t�I?*.�0pv �om�03S��������僵���#��-��E6
���d?�Pm$��)�u��7���9�#��j
�� L8vR�����K������b��SȰ���8��Db+<R�o��2�\[����r:Wc����t��
�&@F�ׁ��k�rY�(����5Qe����'W'� �8��'����+�I#�)��'�n��;;�8��/�B�@���[R.X��l��@?YƭI������m��(��/��$'yfy�_yG��4yznwh�~����<����G�"A:�.\�����(�� �ʌ��AN�4��4�嶺l���@j3� �:B�\������3ޕ=��$f�����l��j�u<�I�F��}�M��F�6�2���v����q����Ƹ�����r��7���yt���y���xR;�g\��T��X)&Dg."���W�4@�D���^���qQ�l�#"}�[4I8[�*�����С3��V�%��=R�\�6��]��<��t��u���&5�\g3�ޗ�K2t'q��杞�R�|k���~y����A�+F|����}ȴ������!ZGm��P��ۆ�r�>)A�u�oX.�@
b���H�"�W%����B�\'��zc���HӰ�q�JO��y���Lq1�����h�ԥ�<] �۪�e������xLu���F�Ry�>�y���0u��,�d����>��s�ܱQm��0�,5z�}�W]7�vP�+ҥ�裹�/G+��oBI��`2 X�RE�ؼI(����ޙ���9��q�aY��4������SיHض9���Ⱥn��p?̍�b�$~�d[s(�� j� ��"����ي��!�P g��Gub6v�ly���+4���ڰӜ���Յ���c_j�	��D-���r��՞�]��ХH�+���a�D��E�%�J��	�:2�7M�Rx�Z��]~,Ơ-)�:�g�r��I_�F���="����	@r/��$�d|��=������������g�g�m=��qq+�x���\�y��S��3��Aߦ�=�'c��O1���P��8�t����G��%--�Rh^VB���^(��Z�t���çd���(�0�߼�D8��_�"J��X��fQN��NIe�^F&21���?�>�́a���^6�sg/������Ğ�ԫqx�z�����ދDI���:
�OH���Ë���WǊkE�W�&S��U�h*�7p�Ea���)��^J�� %��`5Iܐ�'���D����]�ܯ�p�%�s�05�#�}iW{z3l'�X����0g��ۣ��_��􈾕x��ث�N�R;

w�'9N�2��O���傚��� �׹\601e��4/��5�UP",��sކ dL�w�Kg�� r����x���x�����c�D�Zh���¿!�ɂ��\V���G����8�lG@o=���C(ZU�Hz3���o��Ƒ�Z��m��H�+H���WF��L$\���:b�by�����fƄ�?$gM���MH�L>�.mYR�0�%�?$^4�^*Ż=���mTĭ?�����ČԦ/H��bj;4�ْ����b&CGl-(Ry�����2PkgL���4�J�k�$��͹PpS�9���W��CT�����*'i'&'%�J�p�ܫ�Kحm�k?ʻ 	M�=C���ÊM[�W�`��ER�+V�կ�����c��u��,�9��-qin��Պ�\�63�r�7�j!��p���,�#J��ҭ}����W�W<C��"R\M�CNؠ��n���Й��ڀ�a���)��W��p��xr��#!�T7Xݿ��r���m�"1��y���2�<�SVo�ݒ�u{TH�G
��.��-��Es,����w�oZ��OeZ�騸�%��ZJ����j7��?�/��HPQ��`��M�`lj��RߎҗV��`����I��'乶,����J�R�Xk��h
��P������IV��u�6ֳ����o��D�h� �O0�ME1O��@��㈙�,��KT��3�Z��GY��R Je�R�A�v�ܴ]_3I킔� � M�M��Y�㤋b��B3z���w�%G�}��*�<��w0����������[�6�uv���6_���+F�@J�1Y�ٱ�p�&����:s��L���ŇO^{�?~ʱ��Yo~��fTI	�_���%�r\P��o��vD��M/� ���D�����g����',!F�q����"P�J�Ll�T���*5�t0�4�N��.K����kbU��^*���e�����H�/�'(�ǳ�ɐc�H���x�s�~yk*�L������.+�{$��Y��Y���3���y1�7D?8��b���y��<�V��6S�dǳ��gh��!O/�&x&���寚1��H�������'������hG�o�v�ۜ8K�ܾ�[��H^ԣ8��9˭�M���7
[�ra���������}���R�ѣ�i����{'W� ~��� y�{���rJ�8<�dacv�3!�4 ���b�e��A_��2��F����l�E+��g���y�n�dFI3g�遀tJ�1��dO�IDL��K1�.���4e	��`7j��RK�LM� �Q?3	,)j�C�����Py�0*�Qp"^��uǙ.N$�K�a4-H�t#�̜]p�;���7����,��ڤA�GY����2�����u}}��[���[-<M4w�?�V�9��Am���(Tuʀ��K�B�=�.���X��6댍�����od���$�l��j�t���$ 㹁�9���"���Sk+�����~I�T[/A�<�zE�u�X�R��L��u��0�h�f2q�8����C��K�KP���_슝���&,a�kX���ٯ��V�X��hy�k��O�[���������1w�f3�̘��4�9�Wz*K�.��H��뺈S�ڍ���W�td��mk;�o�e&\�����uP_�|}�}k~ʽ�Xd�"h 8S'��إ����5]�x��`Z���؁|w�o���M�z�㛄���}?�� ��(�Ҷ+��:2����bƚ�@����^ ��O����\�K<��VH�E�M<�@��\F�Fߕ֋VX�KSf�x�d�'��5ȭ��Y1�STO��Y�/��捡��k�@o�W(��SV��f� ��g)	��K������
@���^��&�����i��֌`��z�M�;�Y�8n��,�A���+oo�b3�9��D(�́;�J�=D+e��癮��Q�3���t�	�����9	wmoR���K�h1�F�����*�ĥ��yB-o/$�c���˾�����@*}�"�v��E��W	��{G�|%.
x�g��OU��4�_=(xK#5�gM8}��/8+��j)��� �<l�Z1�W����$�� �����e�1Uÿ́��ƾl�U�@�Mg�Z���s�.Pƛkˏ��<�B��Go�s��M�O�?_m�PI�}�ܸ>�H�m\���M~��;c:�w �CL�+�����tMV����9X�X��#E�����sȱv������Y4z�� �zy�����mf�tP������Y��\oWjAf�:��VB��F�d$���c�5Q"�����P�ш�-�-� �}�0��?%�FӪ���0�f`!�X���B�?�tt�q�������qd��ȅ2�e s�>F�����wtb/m������0�9�9�U>Y���ۀ�ԓ�]�Ա!���F*�?�R�*�
�����h�͊i�p��{X0%�|�)]�`��c�:���G������S�R����&��BO5y�EG�G�I�<�ϲ�$̙$J��AZ�8�o�Du���-/(���g ��ٽ?��=!Ҽ�*���Q9b�Z׍0�0��\��9\�,3|��*���5->��L��i�����Yb�%}Tt����h�H���+Id�o|��l22S��=N����囶U�|�s�,�n�@\<s�4'.����[wZD¢���5�+���Ҫ��_
�T���9"��Aǚ2n��J��D��/2���D��� ���)� ��SM���1��:6���C�rc���z�w|z���p�>�7��S.���Ƕnbf0�i��rh��y[�0�l&��r����y{��N�*ͩ�>1�3�w�
Ze�������O}0kQ-R�&�qf�ŹqB2��%�����XNL�/i�U��~)�5{��)��*���8*LJu�"�y��.��D�_2l��&?22P0D�T�������+U�?�(��&C@��C_�!�|�r�dt��İƋ��I02�S��O�[�Y''L�nU�=���A1�<۲���C�W��Q����0�@p�kz�2q���97��b8k�g;B]��`�p� � \� ���F]*�!�����}��md�=��y�kE�$I���99����<2A�ZJ7E���l��q��)@����h��6�x�ρ��˗3����~�d'GU�J�����!��Z�qlZJC�D�y�������׃'U�x�2�p&�ӂ�vex<j-:�2�%}��{�n}�hҏ��=a���Lv���4H�x�&'�~�ɜ~�f�=����J�B��ůɖ�2���t��i���r��h��q��>�n���9��.��Em��9}�,����!pfR4��񭖹,uσ�v_\񁎜IS���_����t�P%�~�iKAז1 ��$��]s����h���S\nVP������ i;9�9H|a�e���%�:�Q1�*�������V�%���m���ڍg�uň��[z ���F�"�h� ����:������+�����!a���aRҬ�[l��!�ζ�J˻v��i�Z�)4P=�n;�9�O
��o݉�t_
9��-\�X������T�T��M�<k|�t��~3jY2R�|)'|��y�x^I�LP�@3A�@����(#���df�kֵ,}C9��,%e��^M�5�p�YlS����[� 1��u��!�����f��j�"���?� yt�ӫ1ڿ8�퀺7�O���=���Y�&��Yy��"��\���/RxX��;�\"61�'�#ݾQ9����0�F�r��U����nSc���UDγG����rɰ��նG��^����Bd�Z��,2�i����(�G��~���Q�����-@�b ��`��6R0�<47SQ� ˉS��/%�J�~�$�r|j�'+t��}Ȇ��Ł8G�����]�>�x�u:�ʑiW#��Qc��.����������a��7�H�����GϬս$k�9ԓ}��'�=�Fۄ� ��Ox�R��9�ͰQj�^�
;��eQ+�;�2Y�˨8Tx�^�T/��Y��|�lD�P��F���6M�^�������Dr&<���Pv6�<Qyl��T��N	"F�\:��z
�+��wF���6ߊ�RBOҌ�g��߼G}r���,0�r�ݟ�XK
��Pg��蜚/JN���=�0�m�ҺL^��[��F���`1ؖc�՗՛���hB�S�ܘK]�A�]*�䒚���e�f ���x�-����H�,�OM3}ߧ�p����
����t�wӨk�!�J�1��Lx����  Hq���ap��t��L��ci�e#���w>OwP���E����v$�r�غ�4��-��~;����c`�|�/�$͜QYOO�{Z��͡[��FV!�ܕ�x����Gj�u�@L��*%�>�w����"������I�Q�4(�Dq�9�rA`K$����L�I�)���n�X��Nþo���S�@����ԭcÁ�R;�n
�KyQ�Ghڠ���:�܎	�<��FA7@�1��i<�r$�r��7 �-K.������-��3���>(�w���n�W	Kp�Koԍ�Ȟ�W��&��m�wP����Iij�$�ƅ���N��oiq�^δ�+�mtz�"%��o���6RW��nfWK��"�g��[8��x2ȍ|i0a��$Ae��<�?�o������[��"�� �� eT0[q}�\�$A�FBB���W���nkhi�K-zgO��niidXgP�T�a����c��#�)�d�t���D�l���?v�����x������d�p\�iE;��%���Q<�9�$V
<0���*��7�*��ň�M���g`�T-�Q�D R��Py��'mf<��5H#5�Sj}��ew���l����^�#���*��
Ԝ��vȽ��F��͚}J�����O"҆)�>��pڴ�����"!�l=��M?��zύ��+�P���ɯ�b,ba���>��xLa�!R�,� �Bv������3
���O�|�p�[��t���iI,�2^W6�BEE�AqA�)�/}۴-��,�n���{�o�X��2�_.�8�	�/���E_�"��j�PQ0J���9m���K�)��(�LEd�t5�P{�������Me�u�R�]����"\��z�����.�{>Cz�*�:'�dA[���\t�df 8�᤻�m(6�����R
驟9"�mKF�E�A
CoNx�dQ7y��Ht��L�N���I��z��hYKrW�)!�Mb Ǣ�]GMSSc�T����X=�UC�뵼�l��Wv	d��p,�9��=P�sl��r 
���??���<5���9pz+�0���EcL��P�+s�n���r0D��U�h�)��8Kf��<�_�UY��z�n٤���Q�C?�b Ɣ$O�g�� T+Ŵ�S����.$�l 4�$��Wpj��n��e���L{����h��������ӐX��X�������	 ^��|(�� 	ɏ�I
�ScC���@|�j������"
J��(1Ϣ��Ⱦ�pŔ�����Py�,�p'�e>d�4*�t����������|��2�r�e�I9�5y��U��Ҡ��N��;-��$����	�]�����OW������T}Y!=O_���eY����?)>l	�z��پD7��?ˍ�n���$<�;����8�p��|&��	���ZY����L͢V3΂������Ή���x���� @��V�;6t�dK���g��2 ����0z ��Q�������Ɂ�'��T�d�%y�ޘ�b�����?�F+J�&2���*�D���c��,�����E�NR?�Q�T
��Kd�Tc�Q��[?.�z�;�9!�e�T4�n�D����&6�iӰ�	�G_���d߈ˉz�սEbM�V��?��$ J�"qP,\ܧ�.h��}�u�I�0��#I����~�݇�.YNt�;���K���4��蛵��=��K?U"��/@C/��O�/���m�0IeF=�i[_
�J�_3��6�.�Jº4^�Tf=�X�ϷÉ��;騻~p����]Z���$W�ݑ���%�~�_�w�#@6�J�4)�銈��ٸ���<>�s��vs�f^»�+��ɱn�4s����Z���`�q���&�.��8�,�rE��m�U���"n�@�#!x3�j2����ՎJ�������n�6��i���yY�!?&�	���^�j�\�C��B� "k:q�}3�f�IC@����޼���'�4S*4|��ȥ5!�"#�jT<�@:[d�t�Ct	�[▩%�R�>j���h�D"���+L'*)�����s��Ӛ�^�v�$��V�\W�O�* �'D;�Pl}���4~wۡl����JQ�Y}�����H��E3�O�����=�x�'�) ���j�v��u�A:	��}�q�s2^���d�����Е.�x%��PH:E��m�žH^"�T���f
X
��q7]��V�ߕ\��h�`Ͽ���!��SM��7��3
 y2�y�-
�R��7^���X�k�\7����B�w<�'��Vj��d	J�mLa��&�j�u/��&9�'����j�z��ŏ��A�Et���Yŏ���T�v���FUzzR0�l���w$��=�0*�~�+w�Z�]����t�#�#�F�_3�r0�!���Mz[����v�8�ɷ��^-:����K)Z�t��>�4r�I�
�d�y~Rrg�^5jxp:_���aK M	v�k��X2�nt����#m�:h42�+�=���V?�����[�P@D��?�s�&eJ4Ⰵ3Ą"Q~O�fĎ�����e�b�P�n�,���[��I�����7��B҃�d�W��@�=�Q�Ǹ���Z����f�[�M���i���O�A����1M�ؿ��U�y=9�x��(,���PzT�F��s�j��Z�	�
��,.�[��Y-B¡��HQ�s���k��V?����QlX���a���/��X�K����?�%H�p��?7b�**�D���I�{"b���#��1,���1��)�܌�ǡ=���0�.���>Uئ�y����yӜ{�y�j[�������x�0Ej�Aa);��6��xA��I�ob^������x�RW��8�|��.��]-`)-W�v���NT��^i�-� )�W���(w�@D4g2ɎJ���A�T�=�9oʵk��
�ʧ��{&'�
x��b(n�B.�6s�dm�O�i,Z>����[����]Nsx�������01Ňe�C���3�Y�Ho��ڑg":��|l���[�k�s"��s��E|ϰ)%!L�`$E�2��@��%���A�^�L��?!/�*�̠�sg��#�G�Ir��3x�E��@Lw��41�º�U�0��j��L�gܞ��G����Rb�b*�~r��^���da�;>3;vǢ?A���*>�FC�lW�-T"w�����d��U��Ǘ��=Z��u��2f�X9Y�w0B2����=�0Ԅ����9O��rL����A��i㨣����)�ړ-+�#�.c�@bn�ҹ�L�YKG�h�ES��Sl���>��ZA$炜�P?��<r16�7P� ԍp9d�Ŵ	Qp%&~@B�����Y�
f
����g�F�wmxx��(_�X~V����4q}�ņ*�:H�
�Ϧ�62��� ���I�U�	���h�-ak��R(#+2��Q�<�x���,�e���;=�O�Z��`��6���lU��'�y �t矗��RFW4� ���J1����2J%�У��?�Zx���"}�t�*�)F�?W��ww��32� �*���B�C|Md�WS�
�{{�5���KliEJ�ݱ
P�ͻ�WrKq�n�������n�߁��8���ֆG����9N�G�#�j�3]b=����?���~��G����=�֠�Ee��NڲeE�^];�Oy���H�/�W'?D�%�V6+�q��r�kI?I�Kn�v0�����A$�PSԦ7��А}��{�0���K)%?�����1���kZ�Ϲ��׬�)$%Kd�D$.9;L����0N�H5�y�+�o~��!Lf�\��?�-6}����fU�-�� �c�/�4��;�}�p�hx(jZ��X��Is�.��v0�����mT3#w\���I����7�[-�z��Kf9�  T9�RUo�� �5�  �S����xc*PB��q���'J�%����g�;�^r�.T-d��eթǅ�`�ۮ�7�W`L1E�Y�f� �K ��2��]Q|����ttQH��W�G'T�'��U��UkH9T�7V��q����v`����[�K�;F�0�0u:�U}ÐSwb,�����Hi��K��`��i��ϑ�[�~j�:���9k��O��YW�	���֖^��4祤��Q�B��ǌ�fR-��/�L��k̰��Ɉ��w��/��4}!�}լ�U��cLǳ�3�K�䡙������Z2��LR�܊x´g��Vb�덠��B�z����O��{q�.ȶ��Y��3�>~p'�p���Q�b� ̉�(/3)��i�*� ��hFE�<sC@YQ.����nvb���'�Pi���o)k�7�5F����Ʋ�k�r;�2������_<خ�6��a$�5��[�{�����	ret����)�W����4#�~|�1�;��:�S�+]�塶��ڊ�tdv�@B�G(�y۽�/�]���xcۮ�ɉG5G�/6&`��+��ܾ�)ސ���B<
y�y�Qvр���\��C3ݱ���) �듼���@�"{�fi��1��{���g���f!����ϵ;����/�TLl��N�ͨ�ŚD���A�##��lCf@4��{-p���u��>�^���}y��Ė���������L�7<m[W���,��I\�����0,~2m�r��,5����&\q�.���ťO�����h���<�����{��օ���0v!�O��̈0&K�2	��㷽"�6�Ň׳i �%û���j�@|<�������Q��PN��:S�����{x�'�c�Uy?s�R0��S��Ͻ��A��"�.��ҧ�N��J\ �b������������h�s�8�l��d����mُN���a���AFƦ,��Z�V�`K[�Ic�&_�@���Y�/���>��$�Z&S����������z�1뜈�$sP]X��}]g����w���0�O/E�ߩ��L,���붷r�}�p�ǪN3��/�I��Y�]�������y�ayz��r�A8�|�4~����2H�]3�� ��|�^��K�項)���}}Ȃ�,�$XI�n7������kl����$�~G�`��]�K��3XzD�8�
����G!��B��,��Iu���I�֒:��P����Y[������B��[�א�hݮ1�y�3��X;��2o���P1�0����,p؄18S��3��~>��pif)I	K��
��'�Y�}މ����L��-�����<���?�P�2�Ru��1�rN,P@�&���{f���J����0��b�#�J�������ڙkU����O��_�Xm�tޖ�	�����
�N^�G�J�7�ʆP_��5���PF�Go�G[��ǎٌ��r�U��1f��/Ψ+Ę�P�v��ul��jK����~F�gO)/G��zyc��ݺ~'�`$Y��4�n��E��(�s/�YX�Q�A��o:wq]�_d��>���!�֟W���*X+�X�Ԍ�J[['2��-�){c�9k�5q[|���h�"	�g/ZfB;�+�w�
���hG+�Մ�>$��	c��>�������I����˩޼Jθ��4r�m7��,�f����:Rv�F�/(�c�E�$m�f�O,=���v'�k+�����9�}(;%JS�дY��)u0�j��{�J,�"
u��c~7����Ė
_c��~z��Mܴ,g�[� ei�#ǉ���/k��mC��cFlw7v�%�gq���![�H��G?��R<g`�)�3{�}�B-a���*I�L)��UbCilF�	����`��!��Ai���ڵ{\]�Ʉ�V�����
$��#�8g*�DkS��)�^պf�k��O>��� `O �<�w�3��@���y��P�4 S�dU��I��)}a��x��P�\��N�b.�=�0�xz Lc��y�E D��:��9O�I��1��>&���pe��$:�d8�LdS��%�����J-,N���9�ɐ��9j��2��ĳ8�lw��F
��
��B�h�1޾�Rd'M��ȀR1q�׿Ӥ�I��k[���WqNSD�rZ_;�kLvi%�g�U���gK�J!��|hE/jS�(:�k*�jnMLщt~��#��o;�p���;4�?x�{��{sw?Ȭ͙��\��{�H��'�c����D�v��>f�C#�p2�c����zGa3�P~a:�QM��r��W��-x�X��
8���4�s��O.]7A�&��=(����-0VI��*r��$�KL�󎝢��_Fz�S�[�Ba@vt�z����5���k9�����2��"�W��	�SnXF��뢫��?~���� ^WVA"�w���3F6�w#�\��V���C�N�乮V|ro@��b2�AG�%�`� ƃ�B� 0���J]S���\�3������Wg���ʷ�t�z"-O�Ri*7]kQE��U%��q/]$w�����jR�ȣn��^�شj����"LW���A�<�޿�P��I�Ѡ��(U��ۏZ�*�e�|��"Q�p�0/,�gM�9ٕ�
�%����2W6����o�Li��P'tǣ����#�C��.xJ'W K���v߻J�=�i����PH?���2�������^�<tt�%�W�Q]8U�������a�(N+V��/}$D���p���p���}G��[�EenkO_�:��*��6���Ϭ;���O`���gLC����� �$͝L��2�)�'��Jη�34r(��QYIZ��F��/W	�'FawÃ���Ѡ��*`�/�Ɓyo�Hso���x<W�r8���~�����ȣy
ߐ(n�ؙ+!]�Z�q��
�����.ձ0s��g�}7k+�X�Q����]*�=V��J}�H-���#^�-�hE����]_�$N��z�ݶp�HL"v�\V'��/<��sA�w��b\ħ����]ެV8�k�0�*n���#F'a�yb�")�� 1Cm�mEZ
��l%��I+#;ii�� �y�#�h��gGy� o�*�-���:qe�
���b��"����Y uA�w��M���(Vo�`Ѿ7DZ�#�����u<<��{OM�B�KH�Y����]�CFL$s�D�)�#�\�$?����p,ie�t/nݾ.�)���
����S��/B �C�Vl�&a)6~��/5oAT���,1��zLm�,���@�<�O�����H�Ԑ�)��|I3�C�o����8�����Jt�A��-Z��3��C�b�P/�M�'��q�O;�>��n��V��=�2�,	*�����Vj cӿ����+ʭc��u�P��S� �F>�LP_D��v���١���E5�T� �6	����ߒ�	3���V�(|D�4s�0^C�� �����ɹ+WJ$�u�R�S˞��\rO �!xx@kZ�J�7��{�D՘{��|���r���
m�6l����NfO���S��&�_npd�Q�NŢ�y�[�.��*+h�~��L�@ �����䉁q:D�a�y�V�졉<���;�䍆��Z���Z?�"�X$����v�;��u��A��c.����v�mn�i�� p��|~I�#*]q�	  Ǩ��*��.D齖�&G���%��A�O�W���x�+D����������P�%�DZ�IA4��ͻ	n�2AӋzW�m�&NqT0��B=�N&5�J�i��=p}ͅ5�|�������u�o^֏īpܟ�1ռ4Z�E��Qċ6�����V�n#ڠ:ˈo�Li��������FfQ�	�E�����}F+�iŉ
�z�>]���(j���\`[葞b���v3�$�5��+��sr
�}-w��k~*�8�����P$&`�B(lmp^U�.z�a��my�yQ��ΡE|a[& ��YL�cdI���JTfE���0������6�u\O�ELFg��ͳ�C5�/0��K[�Y�1s4ZzV���+�Z� -�7��5JgY03�уR|Wï��_�jY!���Hr"Ϋj���\�f�'{O'����01���D�y���?W99�����~&���sd��)���"��{����ۆ��x!�I��lN�)��$e�4{�E1�P`N܂��{�,���i�	�O ��(��:5�Fr��I�
�"�g�˜�>����珪�@v��j�SK�7�!�y���'u�E���9<	G��eo|=(�^���j U.�~j��"�\Mg���Eٰ86����0�:C�c�|����H�5;tM����?����l����np�gV�5"�ꤒj\��-��GX۷�����`�������n������t�תޮ�w��a�ɸ�+��N�:��unvH�Ը����;3�\�+��[ɻ.lI�a)ڹ�)��`���x����x7;�;I�;X�N!�0�\v��!�*��s�Ȝ�
�8��]������^&��DQ���wօ��zL���|��ձl�j_�cԷ^,G��El���˫k+�avG޼_!+"�g�X"B0����3X=԰�tS3��Sh��ASz·2?�ԏ�lK)��?p�S=�|˙���� ��{�n�q��|�r��Y,��HH�i+��-�����)�`6w��v�dx�=\�����\VD���<?��Qc� ='Z��\�;b���v�g���b��J �B�!ۏ�*�ϐ%l	9��%��p���a����MKkv[L(,Y�v�lDn��/��u�~rp�m��b_���&8�d-� �Z�����K��!�E�݆�5jL`6Ǐ�Gp���`צ�H�'�@�q�����d}ZB����ڼ���Y�a�#�t3��GFN��K�r�i"=�^C�=�����k̲7�Ib2��uv�<�`���N�W�Wa��Nk]R'P/W�ӧ����zڂ:�Ž�[�sk� �'r	%Ր��v�P��tj�UP�IH��
6�
Ek�}U�:��c�^p?�s�4ßs��7\��:�Ux��.ы\�J����A�ڹ8=L���3菬,v&qj*}C�O�c��D��a1����:z)�Ȧ@��g"[�E��=�����[x!�������^�d(߲��*�٠����C��D�p<�ָ��C
�y�d�%1��)����D�8	��I�\�
����B��s�gH�[YNDr���o�h�]���F�|D�G�bNZ�"l�F��@��G���(J��(G��J��=��a��L��z'���SWH�]�_�\*dq2<���Z�,^R`�R	��@Ա᳕l���#[ܜM��Ǟ�%*�!l�z~6�9��n��E}H��7L�����˫�6 ��8-��}�+ޡ+���q`��t�LvEB�Q1�ևn��V-̭�KEZ�L�NW���!�^�1�8o-�tE�brm0C��! ":�+i��9�b�2���ENOH2k�!R;���c�|K~l �{/�)<K:��Cᠩ� p^�(8�f`��ͭ�MO	���/Ƴq���o`>�2���74�d�$	��W�����ajO�s#@_�8����������w�%�֬�H���O��b�\��|Ú� н��<�0�Ζm�cz#���=d��kG�J6?J9��(��V�
Td`�\��S7^��@G8�MC���e�(� Gƺz	�~Z6�O�Dz咘Ym��7&��4/2��ǅ㴨����f���v;:�k�j
�o�C�j�z~K�7z���:(X� �#~c��������� � ���Wa� �bȩ<�p�bx ��^�fpm�O�~�tq�yvJ�@%�@�3]�c��؜�#i�[)L��/V�gn�6�9�XS\v�"��arϙA��4mt,,���敐l�Ĝ��"n>)OP9�D���4�w�JF��w���i%=��f����Rs��x�dq�h~��Ec��y�,�x;ߐ ��^G�.����9G���Bx���T7��\A�"� p΂���0�n��޵�����>�~��}�����m��9`�R�D��ʋb_V9�� -��߿9CAU�a�d;��t6r��Y�R��~�㒚5<���{�u��o����6S �:FVw��=��c��6w���ke<X���<�-�L�S{h���>�zr'(�a��OZ�J���S��NF�f�f>{?����ve��Yoku܍�7[#Ғ`#lU��8xN�R�"|
���y��3�P <|w��DZG'�_k𢁬���r$�1G!r8bW$�?u��=`���u~��Bf��^���������i<��2�p_g
��r�A�Z�c��H./�CJ�Է4�($�d_���Ӫ����$�ݝ��ڍܦ���P����0��(2n�հ�<��)%�[w�����c��C�G�I�fF�����pJ|�n�ډ���𤑦�-ڹ��VZK���^P�E(]c��<+mL&�V����o}��,qܿ�1#��9C�z�8��YF��ǚ���Bw��i��0����,��+&�!��?�2�l �s�Tb=��S��$4�t���=�����Q˓<��&�"�"��B�
�)ã#�n=�p�rL�Õ^�9l��rGT����K�|�Fn��Y�D�p[�&��aH��$J�ǚ���<�I�DV~��Ηh㠸O:�
��Ը��j��-iNAnEb*2�6����͒(H�61���~�´,����D����)�2�0� ��ɽ���)� {X�99y���wB�IF$�mH��VdxST���zD��.7Bc䍞OW�����f&	@e֍�r�t�E���� \�Q����44��33r,΅�,�����v6;���;�\�cD.Yr���3�?������é�౫Ӎ|��]�[����b�%{o�iy�+ �8���R0*���>@�RrC*c��K�Q׀8��2�x|C���?��f�-� iW��X�3�B�z�կ�u�ʰ~�&.�$ꗼ%�)�-���-\�j�ȸ�ѓ�mS!�R3�����\��-2��=����
�j;)��=�L{�pxb��C���Yi��c�X��N��q��0ʭQB�q^�|��]��O�"�JB@H��X�L��YƂ�u�h�nچ+m�ն�X9ϡ��0�k(S��'��tM�v�l����ԗ��A�:�=I�t�~�a�xI-��X�c��_6[��9�,b%o�X(�7a�$����or���{�0��t^ ,���0m5}�ߙQ���1{��T4b��?H&;��M��;VP��2��6�-�I� �
<|���� Mi�I|�I@�3�5��A�-m��V������*��W3��U=y�\;]����ӮJ�y�U�0g��F���l����k��!��>2nQ�#�7���з)���/�X���9vFV6��og�1Yo��8dp�<~<�:9 �@�{�<Yq&p�G���ґ�Tؓ���
^��V	��+��֪bk���_�EH����l�	���O
i3�ii�ɠ��l�r������cUԸ]��X��1��a+�Gfa]~���)�_�BcS4d|>�8�揼�=%��D�H�	��*a*B������x���5Z������o���W{�vX"���V��@��x���<|@B�Y�o�.��I�ō�M�Ҽ >�ZD*s���D䓟hr���/����Y(��{�5��I:6�j�\��U�D��M���e�N�f�A�̕�D�Ͻq"���a!���=N���d�X?f~v/Nl��7����F��#x�M%&N@I��!�w����[�����]9���}�Ï��Ќ��o�T�÷x�1�`�!�0,|,g��*�RH䈢�V��5��������
�K2L���e11�������o�Jk�����w�1s��k�b�^>���|!�iICh.u8�g�WE�B��h������K��5um#~)�>���V@��'Yj60����5��/��u���+k;d`8J��F�� �: B��!��B���s��t�69�/���N�ǋι�Cą1��\����:JB{��:εMh��*,�\�g&���w@�]��*�dA�Nwr����N�7B�6������P�� C}8jXl�� �uS!`T�m��w6��跒*�f�a��.�����6��c�Ƕ�\�R]���)�c���.�GAl%�5I�|�ߕ7Ӓ��&bC}��O�v����i����t���^~�Ώ�X��$Vw��k�Gw߶��p���7�Ít�j�a�iQW��IU*Ͻ-���̗tw�S���w�ż)ڝD��"�?� �kH!�z͇�Y]wsP0�%6L���^�Y�,�o�$������o�:�+p��4� *���h�r�
g`j`��)0jî(�[�?�[��'M�]���3�)O%n���H�7�"�����d[C,!d	���C�����_�d.`��z��Ǔ�`���� G郯5��[�>$�1���ݘ����b��K�H5Ժ=VgM���2I����H�<]�),�]�u�F��!r�V�Ƈ�/��	ڂMn�.�� 'C|{7����	!�O�jngC�p22��>��K���0W�%��W�>����)��s�O�r,�لe�^~8\�MN��������꠬~L���h��hWf5q��*tǆ&�d{\��^���ke�Q��LV�e�?Hڥ�u�� 2ߦ��n��b�b������Ǚ��v�,����yq6���_.����栺4�5�h�L�(��˹ʬ��E�)��&<a���#g
�tItH� ��$:�h�&���X)0I�j�,7�ōY�YgN:��D��p�����:����{�n�y:��N��s��.�&j�5�Żt����X'qSV 	�^qˑp��&�s)��i"ԕK:���b��g]��1}i��V�z�?��X.����.�am��(d ���+:7����ME3;[K
t�^9̚=c�R��LCK}X�y��nm�0LT����͆�֗�2=<�L��:>䌸��M"��Oi�[��+�\�P�w�W��Rj[O/�|�L�+���vG�
E��gC��0!���W��e(��m�x��1�E�a��:��WEWI�r�Yr!����]�ou��1��~��[�q7>��`�����:¦)�򃞲�������0~P$3����ĮO���ʡo������y��f\�1�A�����VԮ�$�˃I�N��*jΩ�瓷���",�$�>@g�^K�![0�h��&�B�W����"R�g%Ra���B�M���a�I#��^W� 솷���p�m߁�HA�3���Y�|��$�*��s�u\�E���۽�����5�2+����ǟ(s��R�3��Z��_��JK%/ͩh����"w%��ӂ��8�)�]�K8� <�����RZ�:e�1����)�,)Pۦ���t��uq�f���<�̋c�Xe��]WJ"\���v'�j.I�<v��X�/�����W�6�Z��Т���M�p�c1�W$*Zb�c6�����̨�i�4���D�y�պ�Q�m|Ԗ���w���'A���SV|��)�u��}|�3����C/�T_[G8 -�\W���C�{;4}2j�F�7�;Fz��r�̻��jm]�n�a^�){= �>��~ND�cbQk�C�<�1����ۘ P=]e[�Z��ķ�PG�EjjV�_�2�^2y�'{��U�䯭k��4���|���;VU���S`8ھ�9�{>�-�K�b�_(i�_�6��B�@Vl.bqԎb��&D�4G-N��V�ѷ����UO�n�QQ��ץm!��6��<�^U�a?O�H707A�V���If�>+htu����o�3�K��Һ��7�����$�	�ݜ��2��Z�:Q�w���[`���)��z��u��]�4R�p�n
7'�w�(C�����s��
���RuN��0)�%-/��"���'A���hI��#,��n o�	����I���3��y�0����7�h7�0��o�T�3 N��
)�y�EM;Q����\�#����J������/��BXWΔ2S«i�XZ�����(�:�<Gc�F�<�?�HO�p�?dJex�N^���AODȑ�.Y=��'�����fA�2L�@�]���ZC�q�'��T���NܞdX��*n���l�g�iQaT �+Ӳ'^4�3���ءx�2IK<�hH��a��pɝoސ�j��A#ʒ�N+�:d��0z�(�N���2aH�i�ŝ�83���QTO�l��+��xz��`��/hc����+������N�T��7+M)���Qk&`C�E��z�:[��@R�@4�Z��|�xL��Ư�h����0����K������"��I��R�<,vT�l����?����(��?k4�₢%M�t�K$O���=L�#OW�nL����ٔq"ə>��f-�gi�E:�BB�l�#ɽ�ZE�n��I3�!��b�2K0����m\���)M7��+���wr4��R��6OVu�+��6$8�ޤ�',��C����6>M�f]/_ϵ�-�X����h�o`$�	��Ʒ6�Ѵ�7�gq��Jj�ͣ&�2�F8�Ea?L��1I�ɼ3d�xI����2��M���
<��m�s5�}�P�Upm�[��媂�ҿ͒����f��n
���X���(�+Y��r��G$�:�3A+�T��rqS �y�1[\e�'�ކ�����H�_�Su�*�̮b�NQ�1/�c PX�@�d�s�[{exnM5�p��D�+��c�;��'�\�o���2:��1�j-LF�0f�&�5T�N(.�8�<Hl�Z���\��FԞP�
�ٹN����4�x�����~D��H5� ��J�65��F���F#S:�=o#��H��!�2H؁H��!SpA���Ňƚ�W�ڷb�`�.�R�y_ڮY��EE�����+�3N�BJ�%- �Rxv�b7���*u����䄒�Evn�����s^{t�\8r�Ǥ,���d��(�w�L� ���W��-]��H�Ҡ����+W���`�TRW��nJ�v-�:B2�ҕb����Y|8���O@Q�py�n7-Kn�ظ��3l��Mr��k�5r�9,+UqP(}IE�j5S#?3��B��E��ࢂ�&��8�Z'��*�$x���-�*6����Kӯk�	�C;���oA�:���s�P��nx ����ٴ�o��q��`K��US�G��E� ��əʠ���x�d>�[�GL1���5}���v[�kC50�4�)���,��E|՜�����oԻx�v���w�]�=������l�ጺkEGQ�E�F�����e��%xt����n�"P�_�J�ɺ���w�?R����g�'�Zز�=�ˁ��/�#{s�T�����+옊Cv�*A>�W �ʍ
�Z��6�4�a;�0�B�G��' y�	D��}N_7�V�S���� �Y��4��-l���Tĳ˱��	G�ѦӽW�@��z];���MO�F�4���7��X�t)��w�Iq%8�����~�zz��S�?_���FFo�vư��KP�T����[�INp!4�hͻ�#vPO�_J���7�^L�Ԩl����\�I���}���nXh��k7Ӛ [y?�CY2F5K�ɞ�'@�� C#��WU��R�:�Z���_Z���+n��o���,���]���1��=@e��[Ħ$$�T�H+���rKwJX�E�D�V��ujA�<,��F�*s��m�K��r{YmB�%����%f�)���O�:R����@�a�V����Bh\�I�Qe/�G7n�{s/7%Gi j`E�U^�X��I��ݡ��1�gM���Ԅ���5*����Á���vѾ�2w�a�ɩں���F_����H�u�yk����[�Xoo_1k>�fz�.�Wrh���y�������`7����^�>��$&G���-�|���j���On�l�	7x���4���g9�Fц�e���YdH@�j�S�$�"Đ`��lg��F���A��u�J�ֹ�EC��/�ۻƚ	\���<�\�z�����g?���e��i-��%�c:k���>S�B�]�U��N���7�)�m0ɚh�3ݝ��� �X�-��D8��N�q}�����{f�T��RX�����A��ůBT}"Ҷy���.,�Q<�s�J�|�	>-R'"��� ,`
"�N�'�e��7���>�6$����C��>���Ж+k.f߿��u�)D��-]��R�W��
���3��l�S�T��cFC���!hn�&t�\�v����՚�����}Jy���\x\�Q�w�^Y�1N"��&[<k��t%D�;��E���˴%�/�t b.R��x���\J�J����뙜:�O2�Een�%�;!�_���L���t"�����0���R!lx�a[�Jg�q�8�#Pv�If� ϽNɽs��*b�M�/�	����ı54��Dmn��\ �����`��)j���ZBL(x���E-�j�5Q��B��_�2����wk��<�6+�ҋcf�CQ�>n�f%6.���f�T4D�<�W?����W����\�`��w�]sq�ц��EF�o����]�荦�궆�;��]Z��.ry��7V�@;�11�)Ѐ7R��%�P9��x�9Mh�E�9�S,�^e����f��nIi��꽗����x�¦���+Z	�W��?��@�����'ه�Se:�q��)~�+w�4�$�1��h��P�> � r��p�Њ�mT����,�Ht���.<�n�J<�44D��J���GA����A�_�i�E��DyV[�^	z��j�L�}R��\ߐ�*�jE
,�Lh�����ꕽ́Zu�
�{6�<Jnɪy -��[�%Ǡ�7�f][?MS�м��Mc(��΢�_�����;��]s�pR
��9�ٞ�c�SK0�Y�K?/�-0�*��z�_k��EL��rR	�M �784YxѪ��h�h#�X��$���/�n�A��^<gS� ��ގF�O���2��N��g���xJ��ˏ�!-;\�/��@�gd����x��%�Mba�G�[����6�!���dn|�|�Ak��8#��V�L��
-o��0Alh��^F¡��#�^~��֨
��m�p�Y�.�>=�(�Jd,�����]��x���)��Aꌠ��w����<ڳȪ�E1��u�f	���ȼ�!�ܪ!#D�핚�q�g�0#�uy<�ƸL��
wR�Gl0�&����7�*�Zz	�`�c�v�+7ވ�ksA�r��Ν��K {_�� �۸Ǭ��ɇ�?�*��6zu��X�>�F��~��� �è����O2�Ps5	i�j^ne�|�	g�H���i�����27N�B�9n�a%a��%/gX[��0��	Ք�T%#��g�	۱o7(VP����k�T��x��Ɇ�7x��W��0��1Im�Y�ts`���7v���#m��]x��Z��li;l�w
_�}AM�;%e׼��M��H_�Ro�����ǜpQ����9'gU��»��Zɇ)`�HU�����u�tC��o�H��F&kĭ���X�e�{�����M�0�U��������D�0�%0��6y
�yT樌sg�G�x!ౡ�d�a/�&�aE�#�{��$���m`��f�%���=�3N&W�L�-��O���@�Ƚ�`@3�\� ��S�F*P�f͚<��y�	}!�P���O˥��>e�#M�1����]L�|e?����!X�[�=S<`�(!Z(^�=�Z'b�<���Y��#Cw��/��j�~t$��v��m΀����Y����mz�R�`�����NVn]0�9^\�k��+�G��������0�U��c�=v����]!�������ot�=���K��(.8!s$2�,��>O�\�������B�9���؄eH��<��o�g�#}?�;��O�8Mm��,�TQ@�ȝ"���rnXc�WU�Q��\pb�B��Hl������pH�99� �ߣ1��	زq�h	��`�ޒ�+"Ȑs-Q�����a&"g%�<����γ�q��tZG'�g @zG�"��K�ݻ��qA!	�J�N�I�&a���j���V�[r��R a'B:9�E���(�w�g��U���U�	��n~	�<�!}��\BP�'=| ~��DM��8���r��*��D�ƹ��Ƶ��eX�U�=={|*�7xJ�κ��"=��0�BD�eZ��F��E��T1*g���w�FY0�(֑5)�����	\��)�c롐�5HP���=�)�W���
���$��3�R���-�*�L�7�a�4�-~ܛ��]PZ�m䀛.�.yu�OD#ub�l�`�����j�rU��7d)y��Қ��&=J�Ձ��~7wzr�2
'' f�ʑ��=��L��ݰ�GC	�o�v$M&�Gs����J|���z=L��9�$��f,��34#D�I95}Rn����{�ߠ{4��j���8���)�R��kZzօ�tK�,�=6��t��$�0�	 ��K�C)3M��}y#�����t��R?0p����>�Fy@����a�U���3u��|�Gg�s���9���K��R,$!+5�iW�K���0`m!����}^���g{�S�+��Ѹ�ȣլ1l6���Z�� ��tJ�Ɉ�ǖ���}��*ǋن�����^  �Qpn�%"��ӠX�@e��o���]�P��@p��(<�	��h)uE�_�f�I׫Jӄk��'��ׇ��)7r�T#����:w��#R�6�_�Oj���ghP�'ƿ�#�v�����]���#YZ,(*ao��5�}D����9�0�۪�5�=u�g�F��j"4P8�	�뗦XH��
֖֗Ay�k���p��t����6��:�.Ι�r���Ks�x����}S�� R�Ƨ�n���W���Y[D���Ͻ�I�6U�ތ�?�f���U)o$���*�]@mg'�x�"f�@վ���ZE(�zr���	2j�`g��*��@b��B؃�����+�4d���X��R�Ι��;�Ȋm�A�,�r^M�fW��EK&�E�BΑ����=�`4^� ML���k�0���i��Mz���%K���NT��Sl����A���{�G����Ǜ�&-x	����Ц����C��<��@�sE�X!R#A��ȡ/`}5����#N�Q�Qj��E\Z/��kk���"��z(����&y����� ��;�=鳓���c;`����_S�=����6�����ĵ���	�d���Ee�8��E�%Dt۪��I{�c5:�`0!�^В�v=��A�qx=f�f�����8�h 7�������ΉL�Si<��%�U	؝���c(9ӝ���&ߝ�L @��4�6�y�{�i � ���T�z��&��.г�t�����>ڢ���� ��>ty��AA�cVUdmC�Ǚ�k{���x��'"k9��D��" �Ez�Ҡk���U�|��ˤǵL��GUX�O%�����.��q䓀=<�o^d��Y
���9�b:�ށt���l6ة�ې�;�W�aqv��$����D�za���s��?��4�}J�Y��y<����7�V�љ2	���-ǻcTr�O�fX��E��^�?@�:l����PɡU�n�������>�P��]��+㬒���w�Oo8��H䆿5�CY�~q>�G!��V�<�BC����$5�B��w�.�]��ʫ�L](�G�1"U��ğ�Fz��b��Ν�>k��Eb ����g��w�g����!.��r���h��J"��n �j�)e��{��΢�$�GTpd�Rz�w\t��Fi�rkX�}�ȏ��a���K�ȻW#$Fe��F OVU|�cu\<�nO>�ô�o2v^�$;�X�$����;���=��1����gq��R .%�|���b�U�f�݌����� ���'a�M&�*]o>�.�g��=��t2 pn�I�H�R��1�Ӧ��܈��􋀏�/�g����}�j/��U{���l��� ����C�=<n6J�VA����ʓf��gı>Ya�MB
�o6֜�C��f�D.��2�ԉarB]r34�ZƐ�$ G��*����9��
aO �Cmu��E���Y�Ei�Xe���B=���[�I0��mh����uf��>a��l�6E$��:^z1��▒���8M|3�}��/�Ke���[^	w���<bY��*�C![�$�k��� �b�fϿ��"��tS��*�̫/|dj9�I�X�9(q����"/WО���^�'��o���9�e�ϯk� h���Ě��,m���;�*:4�i��������s��B%8Gv
���v�_��i9Щ�c����W�á���b�$s�T&�U:#���Y��(�����BȼmL3�ٶ�;����l�����_�6�`��$A|��	�D"tk,3,h�3��vr}�n]�֎��/��i�o��f�W���dѦ��1�fPĢ%��}�@\����a�ϳVV1��WR���#������������e	&Ʉ($��V��������=HX����B����4f�>�o� �7F�upyI���r�q�q�KA~����af�Y>��GS��V^ૢ��w��ւ-���0j�,�fw��鴝��P�ۦ-�&��vZ�a�h`y�o����JD��h��-��
�C����c
;�}�����7*���֨�g�no�7�����L�L��9�`\�ǻ,S�� ���r�E�a��Ia�Q�
R�Q����h�)R�}���]�xq��J�Ԃ��	U�n�x����m$�Q{��58�e�ڤ*&��y=�,h����Y��J��~G��N �}y�tWst���E�v&��L����}�v�!3��:�s�3�w�1����t�\�Z�c:>�70�Z����u�3��q�w!ˏ"�bZ�H�gX��ѱ�7\�u)�7�7�-��e1h���¢S��d-'��j�p�>���xv�z]�������yI��FCew7aG�@>[�dW�E��m�0���Ꮝ���e9�&����O��	|~&ϼ�K]
���׷�6��J�Q4�K�v�a�~�|�<TD/v`�0�.�X(��5>�c|Ҩ��`�BnAQ�kN�mhʪ���F�{Zq����_���l?򂕽\�	����Q��/�{��4��=�xC@���lI���wߔf\ԧh;K�H_����)���4޲풦������jK�.�*��L�2�c�ɕ��A�o�W6��6Um�l�Gs����
�n"��-UA �$�\�~�����;�U* PE|m��w��Pc��&N���A��t�*�k�@oUB�2t�c���sZ�C��/��˜RKt���_��}ԧb�{u�'(� �ŕ�m�1��I,�ō�x�Y&^@�3���8
Ɯ.�����Q�D�{!��F� ?�z�⅒���0RA�j+9��^}],QX6�(�%�p�X����+��҄���_��H�z��X�ɒQ����	�w���$�M�K]{�Jb9���S4�
E;�9�#g��н���?Mu5v�#z�-��C�[d��&>ڴb}ԫƋ{�T.~mĐrAu���Y��ֿ�����0�W�ӥM� .E�ѐ
������{k�y(r7��\��B|�o´��t)����q�J/X���x�׻�e�g��Nk����$z����d . ��W�'�K���q�#���*O!�����e���K��hx~�T#Y#�5�T��f��nć����~���n�rw�
Kr���p���{}:��HC�Hx!X��$�鎉�u�L"{��v��U{Ѡ�-�_Z��K�{��Y;�r�6��-U~	r����,�ak�L��K�\��[yPB��X��V\��l��aIU�C�&��Ì,/��*
 x�ZZʬ�^윎{|ԣ4utN �H7\�x�'\��4��xN��k�ل�9�v؁b��,��� ��z��Lϴ�y���ه����V��m8Њ����L�A3�ۊ�����eN8��4m�;�{�wmY��N��G �M�����5o�����%�e�(�4����z���s�[������ڷ�
�MN��bP.�컼g��|�{�Rg�7�0��#뵑�����6u!�~���u\��4wH�Oq�~��E�?w�V(f��l���P8��<��u�7�r:�T�-��b;vh#��X<���X��͌�L�Mu!:'�ֵ���
�p��i����ۧ��������f~��;#�%"�g�z^�|�\X��Q�UGPf��d�\��LGy�1�LF�x[�
א/Y77�}�ܘʸ������*w��h�Y���G�ʣ�q�g�oʏ2�F�g�J�p��`ǍAQd���$���h�?xA�6����(Z��uo��膖.U�v�{-�
�ٜ�XN�t��~������k��>��n+��*�h[n�ն���m�fa��TQ���M ۣ|''pOa)��*�����;�����Z��B�m�X4v��oؾ�y��)� [��+,q$E�3c(�.t��WS&�"%�[�6ofp�Ӿ�ֶ����T6A���/ɸRf�o���7�5U>�>7;�y�{JX�%�@v�I�4Qዿp�,	yTG��c��!ujԠX�^��
�1`���pz����4G}V���rd��鴓�9�fįka��{CA�`����zB�P����,���y]-��U�������8`�]���z步}���!?���8ᰰ���O�E�U�j��8�~��J��%K��n ��]���^DyTρ����{�#2L4pX���o�|l@��F����֊g��H2��1��-/��Ex�ĺ���%fy���z�jC�Ѽ�C���u�e|iH��� Q����X�'P�6,�Iy�᰾��;<#�$�\p����ϮX�����?�� ��0���3��J&F!����)�K �W�Ɲ+;�y����ݨ�c�T��܅�˒_���u��*�y�ֿ��
�B�4����
'^{c63ȅ�<�������SJpM�:nV���s:f�{���f��A�+����:��&y��K�0���B���ɶPDkF�v��qE��dk$�)k��9���{��y=��S����i	�Pg[���,-E	9g���fr�.L^�D�盨2��Q�٫�fҠ���U'�H��E0�>#Àc�n,jm}�n}�Z ������ n�E���'Q;�;0'�'��۾���P_D<ň�N3K2�9��� ��W@����c�!`��|A�1� Ko᝸��;�"���y�<c�d�Ҋ�x0/��<��t5,���Ub�S��|�tJ�n���_q�?U�^�l�V�b�b(�ǭZE�)![�I��zG1-"pZ�f[]�N,�~˰�[XzDIY��:ŧݏ�����F���jR��M_vq>��foP؇��϶�����~��I��<��ɟ����!�uR�y%��(����h���lm��+��nH�E'ߘ�g����?nÇ,0d�=+�|��'l'ި�o�S�x����!��@ 3�3�G��M��w6��W���\��E��b���)�^h�"��,bW�D���}����Ҿ�2��Z_OzӨ)�C�UiKK��P(V�Q6�+�U�e����C�[�r4�zNs�2�J�`Na��z����3zI�U�[��xD�^@���Tf!���$�T�,lV~K�ڮζ8`j����ͬ���|<�BC�D�AD@>���͵����
�w�[�Y0EX�#I��/o8�l��\f� l��\ɹ@��������Ȱ����k���Ş0�4���o�3C`}L��1ҜT�W�/��ԄY�PT�GkA��a�Z[���t�~#5�Ո&�0K�9��6�rې�wo�B��t�q�B�������JR'��$�{2�<%�[�&<��DBz�7�-5���x�Rps���YT퓧ϔvQ$�gT(�8fl�H��E*n � "��iڕ��7c��B�;m�u(�%�)��yB��9��y棙�4X�z��P�qXpj��+)�1ͩ�As��v�������fo܍�}�_��O�}��:q�[tA֐g� vy5���� �;~����d���_�m|��h�(0�S���d�.qc[����=t$z�}����\)y�e�]
�]#{��9#(�i,X&A�}�K~�����v��f�!���T��_ϋcgJ�l�B4�r�v=#�Q�'����w��#�7;v�1�;4"��ܡ%Tb�v3�/}>8%��2��+����o�I�U�B�G9�Vt��1���j18����������\NJ`��f��X�v�x�@�;cޒ��s�F9ew������KtP��-�F1�*-�g8�p���_(a�#5����
�\��ui�ڷ�~�>רFL/�>��Ss5l�w�SQ:�z	�W�d�6~־C�>Ɲ�W���)���=u]�D4��i��3��4^��Dy� iz�;���q/(����F pՄM��-��w:U @랳F��܈��v���%(��G)bi"��4
�Z�&W�3�|�k�X�@}�UTlԣ� �ܯ��@����@kb�%�%�fVo�ƃ�����/?�;�V��c�M��Aш����s����5ƺ�R�2Ȳk�A�.���@�%P�^1�?��K�?еſ����4�3�>K���թ�ئ�?��ä#�P`$T�_T�M
�,�x����D���޽���Nr��$@FSq���+�b��)�^w�3u��E���o=E�_��ai���F�	#&��A��Z$|f8J���]��=��ʀ��7���`�R(��Ąm-��V)Q�&�_S��9�}K��8h�E3t�	!I�qL%���)vr$�܏�'�Pc��4QwY��T�I��E�^�#����X7^�(H_%�Yw�O�v+�i�:�r+n�W7��_@CՕ�Ly�;��2�s�]YϭC�K_�mf���@E��e< �|7'���D~���	=K�4����U9��ѕi��.�0�����E�x�\�M�'(K'�v}�1��cT[�<؜�²;�[�����>��AS!bK�Dc�{������/���dP�b4�]�r�_����B�3�P�l2�qRn��H�e��[g,� 7�o4s�4�~r��Q���pcĂ�(m��K�0#0q���m������~����90�33��c���0]D�9�m���Bk��.{i3���q>���dI	=1dE���n��3�Y�	����ܛ����DF�_:�;�
��$dcz�HxM-��t�Ý0�H
�9H����W����!�U96��-�s�2Nƃ�~2��x�YHK�fO�d�j'ďڸ�M��:��ce|��0��ս��;D���;]Y��j��~@Ektv������A=�0�u)���>�`�$�P�yCB�iJ?��f3�O��oF�G���{M���б�}T�����h�j��`����G��i�m�t�t��f��!�z�����
�|����a�h	U����>�f��2 �����4�����}ܴv�8�H)�k�~w�j��{&c��
USR�h��9Jg����?(�ΐ����х��(^H���1�P�r�r,���b۽=G�?�J�)�Q�w�eQ��AT�ΒD�ֲy�z�b�LC'z���wۣ{jhx4i��7<�#A{�w,�^V�fX ms@�WJ�06�VX���q<��ö��5�<ͼ:	sJ�C�c�ф@�����opF�~|T?�9�R~h��:�F�#���{���({��ga�,v��2^���]w��Q._.�R�3h�U�ϲ������t{�:#m8��[*O�r��܃���� ���MPрW�ӊGR웡9@�4	I�ig���kË+�R���&*�ē��ߙ+}�x�z�f <�%��S�4C���޳4C�J�n�]����Ż��چ��wM��"��R:�xo���N�\��<�}9����|�`Xf�f��M*b9l�޲x_u��Պ�\�Nh��u)
�Ջ��Q�RD҉�EH�����rx�W<�q��� `�{�󦸂 �)�(y.5/Ex���K�z����c7�d���~Wc�xL�ej�T��#�N�V��yg�u��%I/�uc>!�&����$&�:�O�`�@�y�5������o��|�Ɇ{�
��)���1{���+�n_�7��$j�>���I#a���3��7GewoB�4�"��#z{�;	�6P�.~�]
����H��[���j�I1��q����L�N[J��Z+H�ly��q�8��� ���U���^���ôt��ȶ:�=C0��Z2� UP��qgb��_�I���?��TB�-��*G��#�֋���q�����з�)Cԭ��x	�0��3Lk�u=L.QX��հ�IiZQ�u�l�h�Y�B|_�t��Bȷ��T%��u��Р���˦UN���8�2� ��b�G��V��@|��fn�py��vG�]П�ŀ��ZөQ�h��{�R�����ᗻqɇ�(�*3���Ҹe@��������{aF�.��#R�
�\�~��]do �0$�zٸ��r��<����)�����f)�_(�ɉ�+g�j�W���GHJg�Z�\��.�"��=�6�Y�������#W0T�vT;�ξO�I>��]��I�tw^�~�̮DG��|�_�ըl%V8��ō��X8µ�^f)��\��x�(RHxr���?��58�s6�ɽ0�V��N�:�!tɵv9�6��F����n%��̯�k
�)����FF�Ξ�]"�����;��8׫� !E@�=n�55�un���<���9h�X~��#��%N��/nR���f��T��@Xk�{
rz=�H�{S\l��`@���n��bgA�<p�[F�֊���o������E-2��,�]H ��ԾUG@�R�F��/���dX��ۣ��P缒�p(pp�_�!��K�y�P$����-U�1/V��*�Xǳ�=?(+���gA�aBk���V�/�y���P`̅��4Ҝ��/�}2�o�ZB95��]��1q�*� x��+��� �#�?a�y�����({�D�	̟taw��"��3>��J������{L���xZ]��[�"�v]��K6�U3�6���j#�F�4����M>������
w�[�_\�I�4哅��5+�y(��N,6<� �����ov�I�NT���[[bQ2�8�cЦ�zz�¡�-]�_l����r��v��`����Z��KW����`�>��a�������G%;9s�>���?=��y�&�`z�2�:H�͙�>� �@�K">w��.ASl	q#̵��v�J	���u�je�~��Q	��@�ږ��5�D�繝>�5t��VS���̴�����bɘI�T|�����}H�{�^���[5*ք����7���͢W��.$��^�� ((��Q7I�i1R �S �sF��	�K
�W��� Շ�Ԇ�w/�c/�f�DRfp��j$)��Q��7E*��Ai�ƽ ���g���u��d��~7o�3���cL,���-j@�m����j�#/\Xǡ�M!�fQ؀0��:H!��>\{M1�rTfbrmBm���G:�c{��?Z���75bT}�a�ϔ�.��v_ϟJ���tGm�ʥk׊P�vxu�٢Ԣ.Y�Y�Y�w��Kj��n�A��d2���9�^�׸Q�xa��iq�X���d���筤:��T�n����ߙ"�K�#v:aBW{�&�	�h�~u�+�1w��7�5?�#2Y�vk�"��XN^S��'�v+W/�y>=d ęy���TF0tys�@��0}1�[��ܸa�����P�}![�Ϭ�
�Y2���B���H�'MNW]�%�M>�B^d��� �_��0uRXx����P:+���'�����@�5���2G�H)LDl��@RbB����fl�l&�ȕ�l�����%���|�k$;u�ߠt��J�7�6�t���m`A��9,Ф�}����&$yJ#�;��ޅ,�Y R�2���ș�4��l�*��;��$omm��e�̂����M�Ǝ�T�l�C 6�`���,�(�7+v_���3����(̟����&����-[:w�0���-r��Qww(�38'�:k��˟9Sf����c�[/=��D;G_�G��s�ș���˯�n����SuEU�(�hzv�H��_m:�X����;�)�b1��� #�nJ�*]��-��Kۂ��
���y|<l5�^>`�d;u#��;�$���ydlM���{L�Нԭ�ƭ��1ɓ
��g�� ԉ������;%��Jp��u!��ĭ��Zҧ��������X��(uy�]��[`�>y/�ר5y0��l�v�qs�)�W��,���I8
�_@T���jycԄ���p�05���6�U�*1| ܄�o��_Q��}�:���R3�,9٦~:'c��f�������<K��Kei�l{�!n�����@�x`\;���X!nm���U2�WX�]���T���zƍ���p�}�����U�r�14�d�l.)�������$�g��Ha��>@�_�1��R�\�]��/B�i�Q�S�ή�?W<1W<���j�>3'�5ĥ�|�Bz�S6��ΣUHj�գ ����ӊ!Fb�Yٻ�ԛ+b�߾~�t�:	��|�̖"���ٹ@�^#M�0�*fT��F�����Ӣ�n<��ڵW^	E	�%�o�q`{��K�v;[u�R��w�KC��u�.J��mJ��}��2��h�冧O�ODL�i�ZP�[���lt��J7�A��$j}ql��ͬl��H�3�&+��L���j�*��>0Lq�љ[f��]EIr�RA����F�g�z�jJ?��q�Jt����������f��|]p����(2��{���%v[�_��`���C�7��Z9�c����3���'�'�=�=�M71�	��bfc���]kCsr|?��c��s\�������������_Qļ��>�a2i�y�!Kw�����.�[���t�p�tܶ��LW�6�C��b�"�,�6]<�9�U)��q�RZ��D���d�k#��!*�H�CC�/
��z��Mcٍ8Gc��������B�x���oH�����mX���<���n�l�Ĩ�����K���10����#w�2!>��Y����0\�zf���4��E���+��} ��	I�J���M����3��7-���bS����$�����j�9��p�A��h��[Ѩ9�ͮ�G�ex��~�D�S�˟!&�v�x���`�A]/*<n)���Pep�U�>���uL�|�dΫ���2����re�D���&��)�E�[�Wa!��M���1�����1/��xb$H��l���lڶ2NV���nk<^�����Q�� jm>ړ�Ѩ<i��ސ�Gk�T}�����Y��wCmkw���D�U����^��F���~%�8�!��Zْ�`8ޤ� u�i�]�[d�������Y�Ce�|��nJ��	�}�٧���.�0t�B�Qv��8��F������}��R)?�<��Gv?���@�|��D�Y�.��3�Q�l,���������v(����`�䥎 :�4씐>l%�]4��L��-kЮ�5�d���)���;��Tۓ�Ɍ��3�`xM�	����� w�Q~8w�Xϐ�d"C� �-�]������m��l�p3�G�S���!3��p+�z����<~'�VʇNs���*c���}ǲ#k ��ͤ`�5{&d��8�l�U��ж�}g����4��:�7���V�&���MD��l$���r�[]RМx���K�?���<zd���̪��%nZSD״CyPp��A�sw���m�g6�gj�Um.84|�y.�L��~����y��/�����9�`y�@e�-��OaG�^���#�X/�∌b�;�]3
K$�l�`Y�%��n���5���a�Sq�G�|��c�Dg%��ؚ�ct���*ѰtB�G�!���H�U놜o8I�n�R������J���,�c�(�o��q� sDp���p";��T���cwwC��p�:[�~�nB�,r�"�~$ĸ�Ah��Er(;�S'�=3�N� ��0K��G;�P?"�oc�A,Tb��dA�Nw��'P��j��Ko�Z����Y��n$݋7�'*���:a1;; ��4�х�Wq.�|�]t�XS��'��e)����a܅$(4+'D@y�ܥ�+*��,�c.��>���P+B��x��C�l��`Yѷص3\���՛%~�&و�����4�dX����gXVt�F��\�br*ض��W��ɬ���c(zH�F�a���N$/q��aw�L7Obmw��_n� �Ƚ�����~�=ܒ��y�'?Pp��7�~i��d��Yz��������~��W���>��o������A5&^����M�e�ה�C�O�rz#$���y��E�)}�P�f|�����&��U��nj=�=Eδ@�yj�s�AxA�f_,����9�sI�i��=��8tZ��YT��8wIMQ��:{d�҉x;~/ɇ�O��,4�j�%d�S;�Wh��y�<�B>��`��C)��lg�M�%u��=!�r�H����dO���H�!�;�s�T��-x�8���g��8h(Ef�s��r}����0=;%n�|_:J��o��|q/sX�ǉ�d�u��[�4���R��Niq3~V�� 8�a�>;#�z&k��]�m`�i���5��S���̀v,�6�@Л}-x��m5����n���_� ��(����9��O��x�����c��DN@��\�2so�5� ��r�VL`�"h��zGH�y��a�v/f
"p�h��<Ћ��F}��x�$���Z�?�gK/�ѿ�o�P���=R�$ �4���.��w��$/�=ѦB�T�`��WL���>x>CDQI�|�%`�	�lD$qv����!}�����ߍ�\���1$�a���� ��?4���-��UO����2Yا'x� ���b���MY_��l�����.����#	�+Q؉��<nQe�5^z�-�ʰ\�-����[��O���t�w���\^ε���A�EpZ}�9�pN��4�d�܎"tG俪'!�60����F��c��D����������E�k6,f�A�Iޝ��j�߳����$���$Q=�碈h������hj������*$FҗH俦!`Y<�7��񡊃[�(��iQA�@��Rmt�f%� h����G�c{H�:dM���b��'?7u��h��$up��`pU���φ��W��4#ˍ�$a��ߏ�Zc�����'?/��Gv��g�Cչzx����H��&	� F��O3S���Qq��{d�rT�VI
U&�w�G���S�b�-�G q���fqd�CZl[��Z�3x���c��?���l�l0���I��=�O9F�e抲���G��?4��;�����[��$�pD@:�3t[���Qu	>+.X���5N^��& ��)�»����u����?���RX���aR��y�Je�n�}n~X}'3c���J�ܦZQ ��(��_������O�֜Dy:E��=ǧ Z�كH�:�[N�^�i��l����Dtc��&�ڠ�F�/�(�)����-�tfrD%�������K5}��UUJ�R��!�T1�_��-�x15�a��=�p��wZ�d����ABp��y��,�ר�ZM��=i�������Ɛ���By��^>"ɷ<�B��sH�Ko�:�pt���~�<�.���4�N�(�k����0c[m��ݜ�T?���KL%�4
4�b��KZ)C]���lV	D��{��(e�E�-�=O�	k�K�	��lq�3�V�nF"�ņwQ��}�KK`���q�e��N�����5E����_��6F	�֞ �&�WBN)���3�XxfP��@\R&�o?d����s!H����΍~{|���U �s�^��\�}E".�w'�ͳ��9Z�\oG:���J�e����?O<{ӡ^��id�l�Q$���6Jd���U���jt���!Λ�<�:�<���(��,��j$��I��r�UD��s�q����?f�2�������	�~��)�����+'��4V���!�[�md�є/M+� #���4vy񫚸r��Lbn;�5��e����,�����Jf��ӌ3?Vr|�6{E�;�4�pV���Ba�����ED���e3S��Ol�Qo)�Y؁Ive��ZYͿ|�����'������a�>���:��hHg��h�#hj���m����;��Cԏ>����N'�n�XH.��`�k2ny�l���3�Z��v���t��4��J_�%HjYm��Nl��z84)�']��рҒ:�v����hanA<��M����9 ����OZ�Z�����J�Q���g�!Y}��l���"�6x�L(D��Z��0�t�H�D�k��B$����N�������V0{`�������B-�<ޕReT��/�Бʻ�{[�v�Y�zW�%�f9C���A�P�<,��'�x6����}3�Hbl���#�(lT�;���Jc�-�qx�83ˤUn��K&��"�+���br�k9�!�YuaX�9#�4��{w�GEo����2Iqw?J�ʭ�q��7�aE/��ˉ	b��p%�����o~�`H�^7�Õ�Z7��"�<���t��Y�<Q�Ol�f��ˆ_�o�L��\n"l^u�5{�v�m�Xyz��.�Ņx�c;_�c�Gs�D����O"�t�Ӹv���4�&Z�@��RTUFav�)Ñ�5cUת0i�:Ɇ�K��ߡ��L�8���i��H֥�?�(��C�_C�Å�^N�������R�k�t�g2�wPb���nn��0�(D���bc��̱�#���H�aE(��j}bRT��Z8�YA9o0o�Εj1d� �f��8�}�%�B���mA3��#h[T�^�V&~Y5RKJq���mj��H�k�ڮ��.��j&Ms���~;PY�Ă?�3�i_�Q�ڼ_���l&*�:��U��8l��(`�ᨭ���Y�u%@6�g_�YW�H���;̒��DcT~v-Y��a���G:����f5�S���h�~CX�p�AP�ܾ����]f���^�8�4s	۞���"'���2������g�-�G�� nj&)��c��.U�;�T����Y��曺�@X��r��@ۅ�.�K�x	.nZ9�3↑RR��x�t��j5��e����1!S#5Q�*�8�������ܨQ�QP���-����7�$���f\'Ƣ����&K9�D�q�||�����P�.-Z����e����&�����Y*GKu�%���:tY���(�^~�A��c$�v%$O�����9��Һb��	�PL�qJ�Q`{9�@=�0ř�>�3�yԊ&��>`�|[l	���9�F^?3P�����֓�:M�2'�� ���+"��nݣ���=�ȩf�:v
�#lPe�\��Vo{¤�06�b����.j; 'Ok�h�6A� j�ױF(���?�swA�A�C8�H��ӈr���U�>�O�/=�E�n��9�u�����*��WD
��2���l{��Ƕ�˧�+��0��^56K�5�"y�U!�w��Z��))�i�?�D;�4�P{E;���y��0��Y�����L�·�����.30"����G�&*F�>?�	6�וJ�.ֱfR�R;�&_h�Ɖ���6���Ù��G&��Y��q�ㅃ����v���cܥGkX��|�+�4�e�֎]�)��2�I_��Z��Yh�K�rԳ�^qmP[�,�����5ĥ��/�	�C���������9`�w�z�׍&1G�ÝB�S\?fV���t\�yk��Ń��ͼdUs.5��I �����`A���"�Q+|}9��I]艪�Y%g22O#B���eK�\u�$"�c$��n_�d�ƛ����&v���$�O�w:�gD5l��M ������3�*bb4��&^)����Q1�Y�{"J�i9��s�����;)�!�����:Lݰ3��=ep�ť�̊N℮�ϴ.}7��-��c���& f?#���_�+5�r�DH���ۨS��^nB9�e:�&��~������]^s�7��@�~��~�Ϝ�d�GW'������S�s9��|K�Y���7(���SaJ�����H�R��VǨE�UK��|��n��B���^k�؋A�J]D��1^/�|��^�����@��M?���_R��@
�n�����2k�ݹ*�HS]Q,/��j��1�L�i�]���8�)!��D�W�uR����ū������#��Tq�/ɷ�wK�o�$#,��X/Y�#yl��`G�(� ϥo��Br�~Y�x��hq��9��U�"��@!4�����H'�M�?T%~[�\�W�U���-�7�۩~w��+��+e���)�.�E~���,:W�L�M���r>9I��oU�鱳7rjZyO-�P'��Z��D�.� ��De����d����pK�V?����#j�"(e��Q`Z�U�z?�f�e�@}�v����ꂶ(�z�s$~�78��������Ѻ��/��Z�ŝa�\r�Ԥ��Ln9+~��9�O����-��0���4�P�I�j���R=�{�Mj�m���CjeԖ�*�e�E]��,C!e����i}X\8�k���D+хܨ��uN���'d.�W�&���_�[���lY�ů�/[7QaTK�=�& �`'k:>��Ky��_@�IYs�y�5��U����N���dC��Su�s��`�RImG#�7���Ε��P^~�P�w��&0���23��#�D��(#&�qHXPb�O�<TLGg���h�pd�l�ǠǴ^*g����(�7I��,h�uOw��6N^��T�2s��l�}�Z�2��]Bl�h��ZcV{SvzU�֏��m��z�R9=Cn���OR��M�%ɢ�'qf�Sԃp��0.X��������߸�uM>�O�gK���z�����TDċi���û�}�]�ݲ�ߗg�4��o�w��F��7;!��g&� K���=��\	��v�t �}�	`�ӝ|z;�}dnj%���ͣ�&�t݇�o����_+y� �Sv%@�Q�V�h.|�Y ����)|�M��l�և,�R ܲ��!`�c�������њ�2�i��������+��9������3��N�9dk��_LE.B�k*n?`����"��Z=.w��l?�A�����
7XC���/� �B��Xq8��+�a�$%m��cQE�_�Of�X��Q,R֥�gc?�i&�dZ������a��S��!���-D��f�G&h����濉Ki#L�M�>�U����7������>���J��%/!�\��di�����,A����k�@Q�.��8��O� r��[j|ɘ� ��s=X�#a;y�6jo���Q��ʳ!��΂|�S/���� ��_��rI�M�e�UH4��0��5�)�"����6���z�>p�;	�jF��-����+�]@`K)\���-�i/���2#wVc���J��O����\��$W��n%�4lU�G�6eCsF(�������⺧�1����ФL�E�&,� �@/�bL,W�+�_��D��B�"���7����0)��_�N�������9t@UZl��n����A�
z&���i��`����gF�=���§ٿ���RԨ���J�����- ������_4���w�Ϲ��R��s85髗H�VGc�S��_�%\T]n��>�8��$Zt	� /�s�I8�ɟR������NTݿpy�@���7&,�[;>ɓ���j���Woo��J:@���r.�>b�_��6�0^�����N��}��9t�G�"@�ɒ`Cǲ�M;��җ��+�M�=��~v�cД3D�~�,�ʽ)XC�<���!��p��]6�BPw���p�����娃}���\�����rGMV4g��O��x̑���G�Kj���2�r��#��X�Qk��\��q��r�X����p���.��=>�I��h7�& A�
=��)�[L�e��Dl;�4�_��b{���9`l��⊴*��;	�K	��-�ɹG����!)�AG��{}��O���.��P>H��U��c�gj��(�X�X�+	��������?ވ��]���@1���Ol�R0h�VA��}j�����n5��G�>�F���xJd���l*�r����|؋����	��BQ#+�[ Бs����t�Bn��4H�Q�%�9���pr�������в�{2�]�f"��D�?��3���jn�kT{�DU���
iJl��g�	i�4����������i��]K��女�q��V�hXj�|)/�-s}V��V����,a5A쿅)���n����	�.��L��c]�Ѩr�2�a�
�MBπ�Тe��m��G��d`t�v�C�B�E���R<�+9<��4������z��Ĝ*-�`�R��9<��[���_3\Xq5���#��p%��:�J������_{�Y�.<�Ff&�0��_a�[Pφ�ܗ�N�����֘�~N�eS�_y8�Z�u��Җ������Y�/��p�C3�����y�d;�#�7��fAUm����r'�h���gw�A������e1+Z���j`2i,�*'�)�(~��~�ޟS�p��y�oHm�jٲR"K�E������?�#$>DB��ػ�
�ok�6\�'�J��g��a�Vk�мb�%�������Ǯ(}u;u�r+6�0��"��Y�I��Q٨f���bx9M���=�;E[��3���@�-|����w�:�f�������Ø��f&�ѿ��U����F�6�R�7��舊����W�8DdFDb���%:�E�f�W!��}
DgOᦊ"��-u	m{�[+1Z��I.���5��@΄���=}�s�P*���a	s���<>(�J�dҭ]���yY�ˬ�W_��)�+?�<���I!y�ו�p��N���\!i�ǝ���	�J�b>��濆j|�z�:��EQ�${�����_�w28ܫhdH�ذv?RSE����R@��Sl[��<jC���j�!�?|����Z�����e�w��� ��Hh�#!�lYOǮ��[�f{��(�"Rµ$,aR�7��vK�4ݑ"��Zr�~o�{I����E$B��I��N�
�(�,��Ld&P���'Y��	�!c����%��UۢU�d����J&����Ox��Ι����㜒�~�.�T�i'Y�вK�N�6�l��v���I�G�/e�$O+�j*���r��C8Q6S�i�s�j/���鳕L��)��K_��)��))R�k�7.Y@"K~Q��0�ށ�G{��j�&��(����,����}������,}�4Ӝ��o���bZ͗��;o&�'�&g֜2!�w*�]2��T�׮��@r���زi�D���[�;�����گs�T%�o%�+��D_�!�u��x-���TT?�Ism6^�1��ﵪ���#�E;f Y�&��|� L��%ׇ��^ܱ�:���?E����g��%�D�5���]�x�K�� �B�qP*ґQeƧ%U
�$9����f<�G$g���G�[+��!�<�eZL�	ͤ+���[\�|��л�y��r0~�V����a��i���� �
����>�����*\�n3�G�6㾬(���g�$��! �~R�"�}�D8�A�|��g-WY�.yѳnT�����*�C
F�li�&�~?�:���c`��Ы�������|�Э���'H�p�^����zD�������s(t/���.��%'���⯥�<�
����˝R+�XDEk(�C65�
�s��$�8�Ce��I��.���&��N/�>���\��<���`T滠3��񂥩q(*ٷ���3i.�FV����<�wƍ�P�7Z0��X��Y:�\���÷m�F|��o�%�yu�h�C�����s	@����B�!��V9L���
�D��B%&;}8.�&(�֪�IA�.��o�K]�Y�����̺�l /vc��ʁ}�F؞�*5�sD��t����^|U�z���Jә�������0�=�.�:���[.)d�((��վ;�j�F+�;J<v�\�+��T�W;�:�!޾�ߖ�p��U4`k����*�b1/����^:�C=��kLAb��a%!P�tz;�Ś�?j���;"k=.n���h���@.$9a�z*l"E��Z"��Z&�f�6�yt�`�6�+� �뀌#�����`��f�Pͨմ�-�;;��QΠ��56�0Q�v��1
�W=�(N	��#[��\Bv�o���L_�<s%��J�%:��kc򻽃��R�3���f�@N{�T������B���1r�Ú�	��S�Bu0�w��`�	���v�}1f\�
�����j���Up�ʋ�c���z��	��pG!�^�5�2�h�ߝ>��1��hl�c�e����x^��ID�A u"��̈�@CWJ.��:UQE��
�;�w�NY�]����o������Ci���bM3�J�7PLJ`'����\��}���HE�[lq+�n#tn��� 	�_`�S.�����O�P1GC_@y�p�
�����E�+H�zV�	s�/��n�Tf��/$�j��x��L�e�0��!-XYa� `{�y���H�e�{� 
�#w��r�2�օ�PՈ��{:o�Nz_�U�sκ�����EL>P� ̀����_�X�5��s���A�Mɾ��^�c��/�B	Ok$,>>W�'D*�h� �� K�2��ld�R}M��V@l�M`���:p��5sӶL�1���9��,~ר����J����� s�VB S�i����i��,u'Vz��9C�����1�4{A�!1���J�Cr\Z'�h��Ǧ!�,d#;v0���P��Fɸ�7��,�U~ܶ��G���P
�B�#J�'����=p���0�@���U�#�.��� '����y�5���$`���X�r��'��H�i6�9&o���'~�>��#�k�Y:ׄ�ь/��h%��3kP��CR��jՎ{NyluM��L��C�
Є��/a��	2,��|���`w*�lxa��%B��Pԡ9����P�	�쩄�`sk��RX�tOe&�#�{d�#�DP_jj:FZ�Q��7VcZ#�Ė N������)�s\�9�#+ϴ�Fw4�bBu5ik�;JW����˒��B*A}g���j�4s;�f\њQ�4�<�#��TVy�wC.���P"@��纽�zŕ��P�0_/�bE�O�v�P)�czM؛	�GՀ��1K�q���wv7��ԥv��!7����6jT>�����U���>�t�;���H�����1���ڥ�)p��9��TC!%o�)k���)��Y;R��k6d�w=چ�H������P�V�t�s��F��̓��S�ۊ�}}Ln�VJ@W�B5����H[S��� �H�ޢ��0��`6O
�d9�W� �a�H̒Ԅ�?�<i�/�!�t����;�M�pq�n>����{�M{�y�$uf�bծ>Y�TvN��^4�p�a�f\���������S�KS[�4�;�r|[��ҏ�"��0|\�d�e�v�9�&G�D9�.�oY�l*�	l3�ʝû3ׄ�/����؏F`����и@��HOwRy��q��R��j�x@�����i����S�)��H��!R�}���7B�g��W��w�U�5�Fd@��W��v:��JZ���4oDw�}�	�F����kzF�A�/�TJ�K�N_V~沀�.�ۉ�)a��%��Ki3�V����I<\�o��)�5G�fס��R�ƆJ�L��;)�<���J3�����@�1�Oj`��f����:R{+�6�o��P��m���He�,���W�A���ɬ'`��,mL ��?�r�!�*3��9��4���F�Qfޡ�e{s�jZ�J`�X0�`�x����	f^�������x��_+h�Jr�?��)�h���'X�{跾��mYB�f��C6a�7�v9��ꩅw������Gj��s��a�ݳG9�43i�72>��W����,����6�V�z�0�!ϷNx/�F\����0<M��Dy�4>.�@�� �o���#����\�
�ۿ�:/;򕸟�ɤ�����K<�2��F��؊��\,�Ϲz������6���t�P�����(U"��)bڋn�L�!�2ֹh���[�=F��Et�����ӏ���W�d����{��U���,�?�$����^�w�,�IoI'���sr�|�qd28���X Z-�MQ�年������g3�Ы��[�`h���<�%����Ħ��w@����ι�����]L�w5.��9�M���&��I��\t��{XFk�����<%�+ ��X�9�r���mV�r@� ��v#�Km@��@ƒ2�3u���^���j�=��C������w��-�5��ө��bzP� V��ID[��<{�b�D��)�"=�v='y�[Dꬬ�(R�I�rߏ7�1iٝ���f�)T@,y;�g3�Ҽ��dNY�Ϙ4J=fI��v.}E�
��`YS�+��_0�ف�0{`1V��5��|m��3�8=
圌 I��t��8��/��|փ�$�J5�Z�F�s@�2"@.=�o?��)=�D�p�,gĤ��L�|������d0��bAQ(��%�U�t��.F�Y���T�ی	���o��YL������ł�Ԏ| w4{[�����\�Cف{6l��Jy����ICoQ"�;B����I�U�'¡h��Q�U����{�9��x�ʾ"����Q>��>қ���v�3�lj�\߬��P�S����S��R)C��;B�w��f�y��a��˙�q7���W��n��3&I�U����s��}�N���n�7 f4�i#�fvUG�@+o���H�i�����Xc���ʦzp�EAt;	N�v��n�-|����ҀKN9��E"�*c�ap(A��"�o�h�d���cl�/�Cs�]l\ek�ԝ}f�kiC{I߻}�HqӜ��ԁ�;Z'q��q�������+�E+��s�~7*�V��!,���qu���mM��/�N��f��Tsu�ŷi��ߦJ|� ����:�9ͮ�������>-B�ǌ�Η١]ym��Z�������3U��!����B�0>�o_���Qd��O$�q#@�����Ó��n�x�ҽ�\�8u>��4ށ6�Ti��HOt���9$��w���|�<*��&��)2�V6r��f��C}�7�)c�����AB^͢Nϴ�`q��M�����^�G:V�A)�`��m�P8u^M���/�qD,�j!u㾫�ҝ�:p�ۜ|�+��'[�ĺ���mƲM?�\�g�U�6��-�P^e�$:ڼ�Z���+�@5e�)�8�R�-�iҩ�R#�t@��v|�ޣ73qD
ޗ7ydX
|#$Hgb�/xy��p=?�w��)~v�A޹�PM 2T�����������a������1�=�����0������qTI���
ġ(OL�[�����hEa�=��v@_zB��_Ψ�|h�=J�'�4� �\Uns��ԗ�=j�U��Qzxe��ł�җĀ�<�^��meO�%:`��p	@� ��`JF�_V�$&�-ϋx��w�?!��$�wt��j���� ������j�·�I.Јh�@�ݽ`Y�eRxWE��c�y��؉�b~���iud����c9L�U�gQ�{�_����.���W��0 ��h2H|�22
�.���׿A��wOJ��e���ɒ���,Q,�aR�M�P9�{����e@O�PY�rԆ]AF�Td�3��X_Z@���$f�ޝ�� ���O��,e�lձ��W�x�g�]d~H;Ԧ�RŚ�C�W�uZ�W���uq����
��^�ҺR���#����\��������U�2��BQ6V����c|G��������zτX3,<?�H�`�Y�)�G:��$��Q9�ǥd���EؖIל;)���ħ����H�+.�H�HM�4Щe�	3�y��^�w��븺Q���Aj\$<�j�]��*�Dc���b{ˉ
X(^�����&؝������P������$c�M��E�<d���p.1�����B�S�Â�f�Xk���'v�,h�4�[u���Y��`�i�y����
?�y��� �D[
o�E���k(9�ö��%M1<��bR�F��T�e$�TgjM�W\��K��r˘h�^�1� ;���0��^"oW�>kغ��t�����yx>k4����&K��"М���A:�t�H�*�@�R�����m��L\C��`T���u�62�uB��.�~��u������u��ԃ�#c����0O�S��cW`������~G�Nr���՜��y<���B�Nޗy�W*���}韲�Ȇ�P(�Xpÿ�d+�S:�y���!����I�A�8��e��	����{���Ѿ��:� 2JO�o�t��� �.$M.�:��tΗy8�[�5Z�ݐ,��$1L9Q�ߕ'b�ۛgd꼣v����TbS[կ*�Q���B�F�?�O��Z�(��[��������X��U4�L��Z��&D�Xt��Р~վ�C��)H@Dlm/�=&N�v�Ϲ�	Xf�5m�4�m�A� ��Aq��s,��M��%F��n~�\/�H,n���&�>�/�/��J^O�)3�����"ɶ��^\kBld��u7���)k<���?��s�n��`�Փӳ�|����E���^���8��qG�U�����\F���t�U̫<��92��GF���[TR�`I�t�?BSs&���e+�?p�ϥ>�>��~��nz�_,9�vl�Y�K�*^wQ�_i�]�V�G���Ϳ���]�ne`�� צ�������0���I�Kgw-�1?�ϐ	��zv.��z#��4�$[R��˯�+��Y	�Qf�B9�\}Y����$�1�w�*�u���
y�DK�ť�i۞;��{�xwKQ1���f��祌���$����؎��x1�n��BJ�'>>��qN��,߸��_����B��A�NR�GuV���qA�"�.	Mv*~d����Ow@��{����6�W~��퀒M�ɖPŸ�M)��;Ø����b,�ps+�L ��t�\��e��E��{ ��["�i��d�&��nW���A�A��.s]ܭek��6��3��:��<�oB! �q�Т�^i#Lڡ�q�)�o��:y�~�2�+A�3�sl���,��$�C�#�Sq�/��IC��F?�{�0���I����vF$7��H��kFZ'�A�PE�aec���u�d�������a����`�ǆ�^��b���x`���"�k6F�t�LED��]$xb�R5y_Ah���$㦗������L�xC-�X�}���g�~�I�fQ�;�Z����z1�����-ŊGP�������4{=�"�P��6���:�j�9c�C���qv@��V��AI��U�Ϟ�8b"0`]��l�Ւ��j�TvL�TG�r)��Z�9�w0�U���΄>���b����U�P=:s�l��@X>�<F�E�TX�>��nx�!�=�@E��k<Y���U�?�=�\ �%A��/�+���&>"r�9!&1<mw.tCo���p��dR��Z�*��~+L3`WrN��̭[R�o��8}��Vwm��h0{��z�͉DjC��Mm��.���0��9Z���̕zx����������b��iD{y�� ����[˥����k.D!�ݿ>�/�.�,�x�a\�\�)��*�R���_���p,IOV��OP��Z9��G#�q�qYuVf���V3�ެFM��D+b�$�|�oiM<џ� ೧dAU�3H��j��+�}Z����g��q� ����$\h	|��bH)�+�n�%ƝsF�i��B�(
�>D���U�i�W-G��a�U�;.
�vŀ��=�fu*O�9*V�M6P�
��-�)��J�p4���Cy�����|��Pj?8ʕ��<I3�iy�����z���;1~r�A���<�_em'��"F��W�c]ï\�ښg�Bq�/�K	G@JOK�"*7	�t�Vѷ]�E�g��:�ې�)���qi�i�^�G\Ȗ�e�!��bI���_k��~�����N7V7�b�P��8d���"�ت�'�J0����'�5Zf����:�2�*JV��� 4�G�GCf2]?�m����-�7��ى�����I���00��L������ã�raXy&�m�[�Iwp�r
%��q@X�v������d��G�+��9)��9�2�k)�M�I���(�x��,b��a>�QJ�X�ٵx�M��-������ �c��H�D�
������q����ǋ��|T#f�q���oS��f�8���K>����qD�{^1��L[,��i�d[�e>~��X_��B��6��#��?kS�)�wN�62�Ȟ؄��0�*�	8�6\jQb�w��S���DJ��Y��k�&gJ׳~s��Иss#�)z�Vc0,����]�L"��9�[��!�C��or%p�y	u��b�2m�ȫ�������g��U��A����y�P7j��$�`�b�L�xO~¤�<de#�NFz^ڦ�=Q��Hh��4q�"��£��h|p�Wz��K�־�ɂ�)���9�\A~_��ʛ-���\~������6�oeǶ�Q��3���%`qH^�
�i"�PD3۴�wE��'ҏ^�� �V�5�"#�凴-���S�1�`=��H���l*�?�F���*\z�˩�����Jg���I;hâ>�׶��Z�WJ���%�{��|�����Z0�t\�TB�1/b@B���
�VG��2N���QJx��t�~Č��D-�����.ąa�Z혾& ��(5��;kec��i�X��Q:Ҏ�f��E�z�@�4؊���ؗ{@k`DKaglVH�BZ�mĴ��e�	���Æ��T��d�~ؗ�H;T͕�с�Zt�����Eޏ����5������q�ˍ1�g	^ul��p��>�5������*>h�ohE,Ti�hc�K�h���B?Q�������1"��a��ɚ��O#����D�Ǘ��]#��)l�T��<��qE�%�0�N��� cz��(%�R+�������\����1_��7KF�p�U̌��j)M��������U��j
�j�ΖRC��9�"�]1z�;����n&2Oq �;7�6�K�e;L�	��َ������qVTܕ@��U�'�Z4����rUS�z���V����D|��?����0���p����S��ͭb{��H�⾋^��Q�Bq����9�v��$s@9�r����a���z�`A��B�N6�!���-@�N��^;��w;rʏǼmK8=���3��~�d>`g����*�ڱӀ�$�;�!%$��l!D֍� ��p#&���ڙ��㒟�&�vT:��Y&�������K� �����.c ʚH�+:i�fd-&BڝA�^��^�8��6{Es��LvͪED �ÛZ�RS������wXјbt.�Љ���6W���ĥ%K ��=��h����v>+�d4���
FO)�Vбw
��}|���:��5*)�����6���+B�F�c�d�K���^���\���vP��0�
%�����ͱR8�C�m���a�3$��^�m^��$�>��W�y-����F����E��}���&��olP摓�p�	#�;|�!����ʩ�����I��J�Um"rbp�pE�)�ϓŧs?�k/YSx^#7x�d:�%���n��j��Λ���Q�K:Lr��U�K�o�*L��~s�jૄ�_�/wL�	,/�kP�-�}l��A?S�8����6�~���B�H�T���F��~�ݫ�� 4�F��:7���D��!�����<�����k,��s����&��ov�7��v2?��wb7��f�y;>����#Q?!T��4�!�?C�p����TI�L��	�X �<�n�!e6�s�3�����4�gZ���>�>��+VF�ɯ>�+��P'�i�v�H#�1)E{��*X�G;!�O����εEz"�,-�MY<�l�a:�غ���6T���x��#���Z;���Ӗ|~
렆[J6��8m�Imz��/�o�������fz���:��V�%�N)�@174䶹;�m�_�ɺ�	Խ�}�-����қ>K?d"?��v��5l���:`�~�엽�K|�R�J��Y��~F!��G�0�t��2}��	�>�0-�S'�_���-���
�rZ�H�T���9�0A�u	ų=;s6ە�H�m��4��Cס�ϙ��D�%꧅�1z������fq��A�{XI���t*������a�?������B8CQ.�� ��U~N��Oc�,��A\��G�$�.���,���]�Je��qE>j�Z��1u��C������{B�k'ƭ��������y;��ZAd� lXJ�F*���&3M�")ɕ'l�##>`y��4�-U�@�e+��Q��6Fv8�[���w0�Im7u�y��Y�R��Gl�C�,ϊ�*��b��(  M��y �ysxYg��w�!q�u�B:����`�X��+?y3����n��Eb�j�K�d�n�f�h���ȵ��f1.r�M�9TqG=�։��Z�
M�&l'м�2\G:Y ���b�<Z9I1�e�UݾU�{���Y�B+��0�,����[��-� ;��\�e�!�.��o��xX�#2pH0�a�?,�(]����%����23�׺QC�y��5�^d�6p(��{mX ���*rj�Ѐu�B2Y��osT@Yf �l}�]ʅ'R���]�!c9_\˥j�>������*D�vZ�ax/Lt5�g��~�G�#ڑ�H��c��H��/�sw��YM�*��?�!/599��O��7�pz��&�nx2��=@y�t��п�ڼ�al��r�ad!��P/,��?e��Mq�o��,����p�MJ�7Q�mE�*p���:�j�J��arm8�W?)���_�3%6 ?Z��������*T��u~���d�C��;�\jQ�kO�Q���>| X^��X��o+����(Ь��+��ZU�U��+��|���J~�Bd��	[ٖ̏l� �	;ӋI�'C��@Q�L�a:S�[��J���^���`��ũ���.z��:��P�����	T��j��l��P�9�FPʞ|��o��\y��I�i��7��z�c��s��~k�#t�"��b�
g-����gO^e�����{ʉ�E���B�䀁�0��~�>����G!x���
�6 "Y��3]�dUxn���[���c][4ݧg�`|oxa\|�T��V�5��%;�P~���`S��=*���K.�o�%?|�B&�������ـ;\ {�h,}Z�Hǯo���vE�b5ش��v����F!�7���#�Y2Fx��k��ho�&���uU{W�HYd_A���E�/��h3�N�L��4:Ar�����nA܂� ����+a���ʲ�%��q �����L��E5q�����+;�?'�6�_/"J	�.��@o��k��s;~VF�7V|֌�ڱj���d=Bh<��J�)"�$.Ǉ�>�Q�{�>Dz�h��qXt�뛘K�/�{�ˀ�����o��,7�;��%	Ro6 "��	]A\q�N�}N�X��L ���O�����iNM���G��9�͒�x�腞�a��{౨d��w�@�U�N�~.,�s�8�<Y�(h8x+�LI�Vًƴ�kztŹ�T{�h �5��R�������%���s����XWq��$@�OSڸ��e�������W�TXZ�CP˓]�4����3��bT>�A;�`p��i2W�|���̶���V%����r���j�,o��;�0"@&\G&�1g܋�=<ɀ�3��!��W��ݒ���e_KƁZhR�I��?`��������߿��m���a��>;���T�H�65����!A6$��ȇ8�j�F��ݓ3Oߌs��"�ud_[�J�Ւ�e��#4	]엹��\�Z�	U�&|���)X�:8����2�P�| Ŋś���*�$��M�D��5W��1E1\˵T.��U�<�S,�ٙ�PN����4ɲ^,�m�A�6{���Ja��I%�Z�[{�����2w�|�(s	����D���4w�X����~��g��b�
��8K�HE���]�^.��ҝኴ�ćǴY�����f���}c�G�;%�g���jû���t���c��(݂[	�I���x����ǥ=��V -Fl#N�c�p��I� �ɒcz0��3(-���e^���FԷk�C�=m�~�Ne�!�R�vm��V�k3)�Org��Q�n�xﾫ5���q&FT�H*�^����Ԟ�[sy���]����%!:�J�=��`'���Ka�!�'�� X�V�w�lO8f(�ax�����'ѵ�}�p��f�@�*q�b���yh*K��������v�h�l!���� R���Z���ɦͽ<E^#)� T��
��^���]���иM�G_�����u�@\���@�;;�NF�,Z����R�㹏��Ґ�4�7���K*i6}��k��oR��^>8.N�Bg��6�Y���U�seˋ*�fv���<.A^��``��W�
��{,X��2z-�z����d��E� �P�~���A��f�l�ʊNEx�Qv�ݪ��u�{��i����BM�9	!)�/k@:�m#<������Π�Cr�y�a���s��Z k���^ĩc3��MV9cB�B�ֽ9�GRJ#�!�7�k�dK�b_��.�P����ou��W�5��_�4�vE�^Qu�`l�6dz�t�ೄ��H�WF��̦@U�Kg�QXa�= !�Vr�%C����J=C)����NԨP+[J�@�P-���JʽH���+�B�d+��c��**�$`j�FS�4�}��|�U�2G��O��
3��J�z�V�{���#7p��g�f�K����R>c$;�n�	��G��<�+Ϥ��^BZ��	\cH�-Iux% G���U�L�\pz�1��ߢxlk��ih<��R�Kf����d7��O�;�����Ȑ�F�BQ���P����<���iYtzGuR~puZg��mO��k���p�b��S�r}U6ڡS(�d�Tw��ň�T��D�i�m��=7}�Ď�^z���je�y�9آi׌��(���Z��M����үhh}��"�8���R%]�dx�H�C��d���ݦ�o9߸Ռ��o�P��Kυ������ɵ�INo+�4����;[;��	��Ǆ����^�D��J(�����a@yA\O|����I�6�����Bn:g;�6���3MM8�-
w-��	�P�Zh�\
;���o���=F���oشS�G\�5J�r�M�ܭ^��s&1�2.>��"dm>k�8˭�79��x،=��#bt,��U��bK���_&���[�y��3lJĿ�ZXݠ+[fD��=1��s���ǅ�
�d y��G<���Ȓ�����U�r�0#�ZE���T��n��.y(N�OӅ�	���;�/\�yV)��<�����p����n<��ȹvLl��(�a�Ԑ:$��a�H�d�$w��oIǒzƱ�_���7y�{��#�w��w[�?L��u혰\�����V��J�Φ^�*e�G���ǀ�Η�D-Vy+곯�m��e�%��9�n��@�#'M��N(G�qX�K0�|��$2���s�w��E�rjM�pWU!IX5�}�����b$MGB25�	rs�����1�[�R���6)�b��x��#���aF��V^�p�k��i$�
 Y����K>�G�':;�N�6||����ql��G�S��o����6?��/���1�4D �7��� cm�F���K7�[�s��D��\
��"mE�5���v�����s;��Ȣ+��V,��'�<*��^	'#ַ$�*m!���ζ�d��c�#a�C���,�IzZ��1��m�{�A���]v"z�w/H����W�?�Qd��Eݚ��?X�qw��T�E��@{�&:EO�V
MS�l:����ꊡ0�8߸����QJ�\�UU*��5
gA�8����H�M��xJ���!	a��L�ܸ���o��tm/�c�8�I�Q�H���ls����0v�ş����!�+J0�P)�e�wwӊe{�EO��],"�W;�����E�u@ö<���V�e���d�{�
1f��n��x�}�����t*� øe-�9��n�	�aҠ�i�\ﳸ����t���{XL��6��#�t  ������٠6�Hv�@V��SM�~�*|���{֪�4��q�v(;�U�;�Mч��t���z��^yd��3��=���r���:�*�:j��Qn: ��f�r�,�ҍ��4�ҳ�[]"I�C����X��hRqK���ٌ��ēkI��Ͽ貖6�.&39��axd����~���h���V�_Kk��d�2�҃S�@��}��oG;l"��vrR�_�ϽB^5u�Wܠ���,�b�lV�_�7,_�y�u�>J�'˂��N�λoI��@Z���� GIGD�e�Ѣ�xJ�Z������k��DC�;�q�弤�biݡ?����jWINU)��r��xb�C����Mm�����"^�ESm��P�ɧ�����B^�e;�O��|��т�W�PT��$;�}�Y}M��ؾ�-�����߳��� ��^k����@����{ꛪ#��q�ǡ�%Fl9��g��씩���ľ\F[F]�[H��1�X(P�ێӚ[�~��y9���K����t�B_�q.yR�pL��-<
�;3)���gX���*H�{���.���M���b���`�R]c�>@��l����vv��Y& �8����]T�q
~&�-4�#|���Ǝ�_o�B�y����jn���B����Au��޷P\��tZ\�`�d����~�>��QE{1bd�����'9�G�A�
K'г�k�3�"œX�j�9N��W<�dM�����6������"kC���� �P<����٫@#px���K�1˚�{�:�{�9)�t`
7���E�1HǶ��_鰨J+{jܝ�|D���B|ߤ�ӯ|nq�"�����Q���2^>IBK���F���1KC�%]i���X����\�}J�"77�n|�"���>�
��eyz�xN�.�C���K⼽�@t�GY�1�N-�4GTFұ�����}!oi��R3�6�"���[Z)�������'�:R�y����%z�OeZԀȌ����십lH����%�P��09��^�����
��7Bڭ:�����q\����lD'P�` &�`䤷��s��pt�x� 8/�"P�z��~e�� 2yh���&�c73Vdt�'��p.BQ�itCec������ ���2�- ���ދ�cO��F��r�4Y.�a%F����E����X�%��B�TV��W#��J�Df�f�E��]�g�-���]/ٔܬ��Q kJ�"�Ďa��E��7K8��_h��a4%�T!�R�Y��n�o������s7��I�c1�`�j�ǔ���S�-V��B������SY
ُa�f�����j�^jP�0FW��kq%�1CzZK����G�8��cō0���0�+�&Q7�$�xH�����3�g�R$��4���4��m��w�d��Z�P��ߪ�b�O�	}�c�K�Z��v(8"��#_�X�8���5���쵖<]�5SP�߉mDk.��y�Ab�դ��iSi�cW�Y����pءB�3�i�ɛ� -��1gof�)�o<˼�낕.ͷ���X�����O�o(-������\2pv�ca��Q=��)�(̌�^���W+�ެ�<��)˙�A�+�ֈ�g���;��h�{��Brk�e�\�������6��3Ps�CM�Q@��R�:�Z��]���YR:��� ���^�U��a�'2�������ǳ�uX�¦��&���8�O��䒁B��|����>>-��XF�fJ'���O����%��be�T�=5K��*6ީ�~������%�&Q�~v�8�kY�p����!�"B6ޕ�@��8T�B���cnm(sP��U�Nb���5�N�A�n\1���#���������Rԍ7��^);����%(�0�ͳ�����]]-8x��-}�fάp�Q���W]@2�.lҡ#}n3ژ�B�C�%�E�;t�64�hoV��,p',�$�9�e��K�2�?K
t�X�i�5vA��j�	�p��e;MO�r$�a⎿ur]�Des3]�r�y�׼��cX���(==Z>�c�${g������#-'���
�M��Q��rr��,\�ǒy�e	��n�3X8�g��e�G���(t�k�A�9M+Z{��(+G���^�8��qsD_�0�#D���0�C��
���v�R����!uzy;�����v���1�S\��I�{3N	��{��3�Ұ$1����!�Q�o��{B��(�����6f��ﻜ�OG�-��8�bz�@Q�)�?'�z��O�Č�݃��@i$���,����Ϧ�F�4�"yI���5�A�����j�:��D�*n=��`���=��i,�y{���RZ[���`|%��	l���|Ų�[0�N�sk�S+��t�Rk�*J��Ht�h+HƳ4�*�xs��\�9�N��W�#]R��J��LĽ�T[�f��-�KD�7E��阷��U�"X�2k���$pt���߃�}������x��.阝ԣt��{��W���	�!�@�1f+y9:&�-��~>]����
�ʧ�����P(̴�Y��=�k�����^=��� lƲ�YG����zܩ�hݣ�����`J*���1���������9�2�0�E���>�u��Y8�pN�~�ee���OoV^"����*�Pj����^R,�Z������5<��v�ӈ�|�r~��/mI�p���E�o��w���B9�_y,�Y�9_~�G���@K��W��gI_�q�u��~�Pg��:���".�)>�d����&P\1��)�^Ǜ�l)�l��n���~�����'�>�6���~*��r���0d���e�&e�ʬ�����|�t���bJ�0�Lj���?z`@G����D��K����$���� ��tG&�����٫D˪��Y��_�A�yZ��ԁ��ـM>܁���j�p�7g�vqB�/���_�p�g��c.�/2_��M�#C�6�|	
i0��쟃9W [ ��v~��#�۹�C�&��Àt��A� ��Lf���zS���i:(C�dJ�. �����<����-���I��d����i�1R����p�p`��U���_	E��zCS��yɩ�̐G���[�'�D[(�ɸdc�tv�R0G�߲�P�F�ŵȸ��\~�p��T)fǜ����.�^�V׍	|�@�g�i�HU�:�ק�\�xщ�㮤x�|cih�l:}�J��ZY���`G�iw��甾P���s�d�u7�?��mZ�T.yd�r�I�6̓2����9Pn9�5)�9W5 T�%*)���c^��ƣ�}����Dy�(��d֌2 �ve�c�z^Ե�K��ǐ��X{��R+oz�xC�]r_�24�6*�W��u���5��C�K�ъ�^ ?7JL c'�l�}>��#���W$g?*oǧ��`�*����ʬ��$��{�d�4�g��-�wR@��}z�����T��<���9���<7�����/?�I<�ZoLn)Uu���4m9�PΡ�
��h]��aF��`1�ā���f/�Li�dcΰF$��������93,&����<��>���GL�q��ŀ���/�[�QwF���w_��Iף̀�a�YZ�?���*ʁUY��^1��K4#��d��?�EK5��4c9��!����?�.�Jלbr�d�j��X�}�>p��7:8!Jz��P�S	2�L�=oK?��6T{~o����V{&_u2��P{#�0���0S����C�Í�Ӊ%5��3�W������K�i�!ng��@wZu�Cj�[<"��?G�����[<��"��<u2�A���]#;�,�/�IbH��ױs��8 �������Z~M����*��I����g��NT.fê�ټ�N�z���˃�Yd|2��<�������)�c�7���Mȥ�ށ��$�f��y}���w1����E$�p^��5p	�������mE�H|V`BH�&X�f��d��f�,Zqw��i���G�P?�(y�9J��"��堜����%�1+�}e1@��9�K/�[��6�د��%#�w�4�����+���ޱp�q���݅�rvl���s&j�{�e8}�^[) (��x8�m�<h�i�ǩ���h��*�\VR�9��˦\Ĥ��^L��?Fy�b��yv�;i��+hq�O�d��s�}Ҽ��SSbz���W�?+Q����X�-�j�*������l
�}Q_#1�ì�F@�e��$ހ�-�C���?�����OϬn"�w��^��h`�2�4�M3���&��Ŗ(?�� ���b��e|=��N-��O�D�~C��ߡ�L��_���~��D5;=N&�S)|���p��I�Bf
ՄJ�-P���|<X��.Vy��)��)yg?����;��gK)<��Һӳ���x�i��4P��)�fǦ�@2ö ͊?B�_����W(࿒y��mS�Ē[�e+����0Oj�?�5���4*a����ɑ�>ӊ#RY�EǸ�_p� Z]p�{�)�F8Ǩ���e֥��_�ʣf�Ҷ� +�ׅ��fڧ����_[! ���+���+MM�p8�!�����=�)�Er�Ɍ�<.�֘��4#^D��g���'�_��-����#�ݨ�� �ǹ�e���p`�p���i�.��R���YS	����Ok�3����ܛQb�1����AH6.�XJ���)눢P��]t���]�A.�ڬ����X6�G�Ɔ����z��� ��y/z�y�V�ͭ_��3Ү��:9T��{�_<���^��J���brYS��/�P�L��y`�C�ؼ���Дh��wz����>�sG��ˢu�#�m/�6>���Bڡ��^�4��tcb�������M��#4x��tF�Ci
{�n@��kd��c�k�z��*{#'3���Mֿ3dq)��W'�Nn�ڈp�x�AP���@��,艄��g�<������l�O(w|��)j��i{q7)�5MឮK���3�R7�ꅾ힯��Yo���XT�;�
G���4��j&V��;������A4��&��d6kF���W�{���MA�Ju�cI�A�a�G6޿�U�2ѣBO�J����k����|�Qr=�N5��/��kȡ�g=~�¸�sh^���\�{!mT���A{�N��k�4.���5�V�}yd�8��E�4s!)g���[�N���z~
e�uMZ��B���N����8�k
$~����4�ձ\���G���
�T�ԓ$;�\�"�"�И�������jI�R�8���2�cn��ߤq%"���~�(�� _I�h�=��T�Z�M��F��.f��vKұ���k\`���z�~��M�ڧ�0�I��Sw�r_�ew�/@����z�:�>z�'���|��)�ܮ��8��ݑ!{�W�4�:�âֆص�&�G�@s\\���@w��YJ�AÚ���-��.��#��� ������Y.�7c��b���^�!�4:�'�g�9>����(��Bpz�(ζ�W�����h��n����%�аF���oV�M�a�~�\~��Q�X�X��S��k��p){�t[r�E&�����W��%CMí7�w���w�!wv4H�#gF>kJ'&hj��#�MǗ�W�7�!@�h2sO���z�*
�Ϻk��c��l"w��Q�z�U�[I��|֯Z>1^G�e6�7o]��~��>g�җ��Łrg�õ� ǐ��Z�����L�є�l��zYr�1�����^��͌��*8��^�(|{΍~q6O/8��#��^�8�;��q#��%3ȸ����_M<�z�>��"j�/� V�WYj&9�{~�:� ɂQ�7a��/m�+p�	A��9�z�����[-b�5�ʢ�>Tq�A5�i�1���3e����Z�'m绥��z������־*$�a�6]�%p}(З����1b�T��E��+ =�ә���SHd.u����T����Zd�a�����I}�6WHZbOn_m�O�H�۫З�g/`��޶
�	qӧ��A��@��7Ox�A�����Q��*`:R�DO`�槎
h6�u��Vm��훤u��/��Wꢤ�8{��Ϋ<�n@l��Tw����d�B��.x�O��v փ��B@��	S�b�p�����=qo�Q��^��@�	}C4��nt�/�K�q�K��P�����u��1-�����H�"vŖs�����X���}��?/��<��M\k��xa��`+EF�*��%s�pk	;ބ����J�٫��Q�m��%i����$�l l�X$���|u5n�D]��̆�oJ����G�5N#]�?�DY@IN*���)4`ksZfLv�&�F�o.�^�8�ɇ�J�,��N�ڸ�
�<H��e�{u?�7���Y�1W�.�'9��T6g�S���f��ţ�J��qR,{Yܳ,���	<�?EY��?<>��z#~3b�S�P
E��IC֕��������+��	x$�;Yr���KO�N�F�
@���k��:��A����?�hx����Ж�� �f���,,�.��`�6�9�S1R�\u��i�G�y�sXr� ����9�f7��f����R&����	'ԉj�k^#/b�6�[N.). c|��E�A� �~¡�D�7(.dF�$M/K�M���آ,����4�2d��-<U7��ԇ�����#h�>-&a7Ix\�G�
u�z� FE����c���S��R^��
���(c�M�7tQ� � �!�dz��}�Ze�
�]���~��?�G}�ó����D�ig��tBTJe���P<�E�1���":d����<�� ̧D��`�쳞�����!t�bOJl�sg2��p��`�cZ좟����!�(�N�sɃ�}mt�CQ=|�B�K{ǩ�����#e'8�D�{�[{	1*�(��eڛ�� ۴���SI�?�A� �&}�Y'b䚭�2�����۴�;�̺#QAXҏ�]Y�S�:-��L
����cC ��x~�emR��^X�T<!�2Bc���V���Q~���V��9g��)�Z�1k+�-��L�격��������C�^���	��T0=��HM���D���u�O/�&xT�rAg,reX�)���,��b�q?�,�����N�d�JO��m�1��Bf�g��8Ue`�����|�6�]�3��gf>�(�6�E3.��Jd��ׄ;���v_��Q 屽�h���%'t�3�7�~d[|�+�A'�@��]˲#=�����L�=/�9Gj�2� ̺��PT_:&�J���tr�����8�n������1���x��{MN;���5}�͗�XIK# �dXi��������[>���E��m��/�4$Tf���}SH�W������;(�3��&@d0^�Iq����*�������w�*�t�K����U�N3.���>�%�U�|V� ^$��C�{�6@,����ly��E��e9[E�{2���}8o	�Ky�&v�x;^��"#j�zQs���P�>�e$��"��yUv���+>�z�#���A�C��d���$X	�4�ֱ|-�j�i�D Vp�{\ݸ���t�R&��/=���'�?U�����l|���A��j����ۮ�����L;��#g]��µ�Aǜ3r%K����y�)07����V�C�FX���?Jw�7ѵ�'SVd|�+��2��\�\\������9wJ�*zPIQzܖ�C	�s�Ƒ����S[��"^yW���7"Q��2���\�)��۹��	*�,��<��r�z���f�����߆�wN2��E�M�л��7�U8�)}#x�^ԁ���=�b��_xV�l�����2l�^�<y���Q���s����cF�˹'���o�����0L������J�W��	Zx�\�%5�|Q�a�G>0�NQx�RC���-�&��`Ӱ��H{s�
ل����:�.�F&��JN�qs0.I>�C��1��vG��ʎ٠$`����S��v�P;`fpʛ=}�hr�
��Ю�TW[$�5�F��r�p�9
���!%���:Wn��2S��(��[X�9�����X�p]�f�Ti�"x9}��σ)����H� d�.���λ�,H+����pĸ�B(UJɣU�}I*Lq�7�6�N/�,�-5��v�$/��Sh�q��,�{����w+� 2>��N�H$���IA�mUM�$�����*�V^Q�GoM Y4F�~�G��[S��+��M6��ҩ{����1�o1ު�����ց�l��z���
���!%4x�^|�Dw��`s2B�[�n="��|�q�m�6���)��M�WQ=]
�7�g�t�vr��ť�o�Cg0�l���rּ�oa��N�/�*�+5�S�%}�RۊS �<1+�e��-����zG�l���ʶ,���Mr���w�8�D�@�]��w�9V:ة�aܨ�7������3*{�4$0>P�|?���A������f6J$U���GS�rY��m�D���a;���-q�ոE��$�b	�s�L�Æ:�&,�rC{�B ]��#��;�!�x���p�j����9�WXP��ç�"]������9�������k��F��o�ϑ+��zpvN�*9���g��zj����R53Э� �ݠ�7'�_I�t�Q��0����$wֶ ��%A�B��'�.����E�7�G�!Ӽ��|�&�@������R��A��Mh��9�8����&N4�(��ٴ*W�R^�Dd�*&��W�Cյ�w��p����*�z�4����t�߿߻0�	)�<����C
s 
U@���zR��mpK�'>�����gF���\���s��0�=�/>��1�=Z'v�W%���ġa9�����%�qS����Vc$�A����l�芟ϱT!�n�U���տI��_�S�3M2� �%�/W�`��ˡ}��G���?	�n4���֨&�g?�	�(��o�6�h��.ֹ�P����+��ĖJ����E_���D�nܴ�Y߲>��%@Vb�	��j����1j�5su\%矕y�����㰅����j\&��g�%_�f� DX_�`�{�A�z]�?�JG�;1�R�1�h1���՗��p�C/��7�Zg��˓	p�%I����WEW��t��lhxc`H�U�/X ���pI���bs
������bn��ɑ�q��;�֘�����o#V��a7�C�}?ʦ�u��4����5/�E�	�(����7f=�x?��C>��"5.7�����`x���VY�VeEi�G��%��Nun��l�EMãƪ����1�����SO"�e�6o��QE��hb�A��5v@��|�<�2��4+?�qf�w���=�ܫ�b9c̚wx5AB+>���M������y��n��Ư��|��ǻ��}��v�qd�6�V��)=��ᚪ=���DP��޾&�O�pr����bR������r����z�J>��!=QP-�[9�5�%Ťe_��_��`���7�6���X��5 M��ʬ�e�}]̀�D:��Nw���A�њ�R��Q��$o�~節;е'NK�ې��W���Fes�5or'�����{Ch{��p�5 �;���7��h*L���D�i��S���y|�opGV�;7ƛ�oHr]`շ1-s�GU{�hY-X�ۅW��L���L~V��kᛷ��TP�,��θ���w��BY�n}�j�8w̉bԼ�L3Y?�c~)�Q$�E�l��
I�����/��Ri�(4��' ����Qw@Q������W��ݝ�ѧǹ{QL�@�ˁc�&��U�������윐_v��R{�b�4{927�u9���s���\��U����~�rmS�����&��͢j��&���tؽz��r���zX��v�F7D�ɒ'h�$��2j_���O��J����?b���A��ǮA�7������%�s%>6���ֺkt���s���N���3�HSdT�����mj��s��U88RP���n |�H���l�,ktȽ�\2Z��n�6�A=��R���v�z��A��s����u
T"z�ԎS��9�1 �� ��rsW�!0c�4�ы�(��j���l���g�׼gMƛ3 O��%j�+]��=߷˳���D�JQ�S%����ZT���� �ـ��I�� ��Ŵ��@`m��L�u��" )��h֓�c��C���(�`���1=5���R/�X@�����"W�|�Z�	�c��FY��-�ː��=�xF����cr'����	S4?j�u:��!fء��C�>#�̉�˾LO�K꧇�+��]l�TY�\��㉿���{�{`�}ʣ_��Y����.��{��6�
q��8�_+R��_�3��V#<W7����.s񤲇l�A1����5�_n�d�D��Io�����?�F�U0���H*t���f=�WI�ݪD��MSO�/���k~��h}U��$��n�j&`�w� W��_��	� 6�U���V2�����t�+{7Z�y�v9ߜ����-�N�r���hݤ6��/ǯ�x�Β���~oh��f�~SkB�W1��j��˝���m��XW�%�*TD�r��)X���]�gW��R���W�1�ܞ��Z�"�����#��б��H�8��V-�2s܇�*���bm�݋�
���\.W2c�4�s-	j$X�D��H+��l�!(l��r�����g�鞆#2=P�,A�P���;+Cʻ��U-�r���5��r$ZyHm�i�e��{ �
�b#>[�vY�V}֗g<�T4 A�����i�����p�]����T�#O��7��c:o5�X��ȢӍ��顜����t���]�Ƅ�6
~�a�DZ���Ӱ�(�ro�R
Νf���.�V��qDP@|�&`M����a�h�O��a^���B7GZ�Ӵi&�g;�b�~�V��a�_��}>ݪ��+��\�nڐy���U�-�{[,s���e�g��{KL*M!ns�̙�Z�udw)/�?���IR���\`�ݦ�ø�r�����cg�^�'_�O^�����}O4���	QJ��5�z~G�ʨ�ѓ`�����2/�Έ�Q$�%�Υb��bt�t��:H!�[���WD6�{��rR�s��i�^�t�ġ����2�L���u�F&�ώklBw�f&�[�$��Hӟ�7��,�r���}/��;��F�V��L�J\Ż�3�2��%����yi�e�Y����W���dBl���b6[�h���WvЌH_�Aܝk�P ��ьњߪV!�<�����,}���g��`��, U9w0�=R�'B����08����M)�̫+�.�e�DR�Ƨ�����4��6�M�D ��Ej���$%;�����8Z����r�������sO��L����7�+[=I˟>�޴������������ڝfS�t�����X��r��	B����Ffw�KO嵟�K��U�Vq�&2�"$�;��I=��EE�}c�LQ#Fy}]h2!�3���}G�am|��?^6�qU�G ��3[��]m���KCm_X���h�z����9�Ѻ�����ܭ���~nC��ʒ�ʒz����~+��N��O�uT]�����bb�r$^/��V8Vs����<(�����vI��~Y@�~�?>�!E��~p �����]�F�X�:�~[J�Q�>������e�;�'Mx�+�޲[���³5/��UIN��3c��'�!Z\yZ��slr�nqv�E���Ő��m-%�J��{�\��U�'B��׫z۱��A��]��A�WIr3�ֹDb�Z7�}������F�H����E��Li���a\�6�?���̋��T`妘�W�ɜ����
p\=*d*mO�� Ѡ�$-����#�>��2�� �һ��&�aȫ��"A�WP*��Q����U��Ś�:���T�6'�?i&Ή���2�:��� Ĉ2s�����P���p��Ш�#lF�/�B�
N��ds�ċa�EHRm3��W�֍�w�2'K��}[��W��p�H�!B�nB�.qB[�=k�偔gv@Z|k��a�%�>�߲"K�DP!�F��n��s����*Ȇ����:�qԑ��V� *�6;��3���ʛ [��,�t��&����S6�+#otɵ��Yw{�Һ#	�
I�d3�:@������w�ӻb8��۶�8�)�wǷZQP����e;0��Vz�	�Y��m���L�ư�}XZ�%s���N���Z����
.�G��^�jj� ;�wo���&Z[��b*�9��2���_.�	����_���Ұ�H��.���YUl��A! S$�զ'QQm����D��X�k31Z"m��0�	@)
?�dd��5.�۳EJԈi{� �?����m�߸��X9�ٴ�nC���<Ԩ&��Гnu�pG	C	�e	@+O P�*$i����f�$n�C�]]s�|�x ��?�FUX%�i�e�D�E Nј(��j�ѱ�����SS���X�c�A�]b�	���K����+I~"
�i��R\���(� �*)�9�K��F�����_�%�����N-�:���|K��/5�X9��q�XE��˻�3e��/�$y���>��EwÌ䪤U0���z��;��C�7��>��VsN��h|�5|��=,���7�X>��[�*����B���{uH�~:�#��-R��6X�� e��&{�b�/7�z��,U����S��H�!�/ 7 ۄF��f�Ӳ�S��a����'6���`v�?��&�ʚ���[wc��jV��.��~~���+N�Y���.�v�N���"DC����N����ҙ��%Ƃ�7>�(Z����%]�::a�@\~J<�#����=�R�-�@^Q���ʂ��E�hq�rr�iʴ�tI��o��D���V>�<��$"Q���Eag��ٮ�n{��6�̳��#�sxW��)Qí�m�[�Л�.獒prq��T%�WO������b�w����F�ހ�� 7O���y�c��e�������=�-q@PP�r|�z�G�-/}�৽�μF�!����/�P4+��֐��U�jl���s��N܍�T(��t��[-�'-�y�/���E��g�����Z��2��;�X��Ϡ��T�K�Cp��87	�7��6+���C|�Eu�����S
X�)c�Ӝ��@�`�.m����VS�TscX�3����)��U/�ͮ���+�2�_,���O`2|��� A*�,��.e]Di�W�ie�w�{�U	���U���<���(l�V�\�O�Z�RQ�'�Ζ3�2V�ݯ�c�zĤ0
�Ɖy��Dɿ��4��H�-d��kgMP�7FGE�=̜���ݳ�M}�7Ԡ���d��Hj�h'E�<T�L!�*#` 	�g�k��II������T�Az�e���7�'xH��NǑwvro�J��u�\m�Q��?�G��Vz���__��׏)yiy��/&ؿP(D���?j��G|h��#��-9�&6Eq�)4�`,��	�n����M��FB���o��qF!wl��t	S�����2x5"�T����բ�7*'>���_�~�+-!ߙ�r��s�6)}+!zue�2�j���\]P�;��n�! �S#�My�#B�J�F:��	�~��o�$^=�7e�H�
�e��n��YO�ƥ�֋�+&����ne�J�,	�T��h ���N@����z`�$�QA�z�>�(�/�)�uI'���/dt=z��ȳ�
-�\e�&y�m]��2ڱ��-ka�[��=A�/T���[uŝv�sQ����~���,�2�!1�Lh�A�����j&��L,�t	#�������?���[�F��0Q�������z
���%����喐'^.ܫ�*�`:��w`�p��HW{�5��yo�J����Rn��/��P�}kNp��(���L�m�	L�v�D�k�1ÂC�xhV�TQ1��u��6�PZ�d/&W��r�3#���i>v6sR�׵�����\��̴���S}�7)T���L�����v���0 �g�s{`�-�K�y�i=	���"�y�,��f�E0ŵ��okVn՝4�3t�OH��O�~r�@2�θ���c%�Ds:�w��s��y<��?�y��'鮸�EUz�ۦ�>���w����v���C앧�#�rh��L��]h��cLȟ�_�~�J�"f^h���P̡N[����U�=�����R�}�V�B33ry�1��E��J=)�K��� �������)(�̈Ю�v�s�/6��}�2{�A�"���H���P����,^���NV:W�{���d>��<�����{��Ğ�'̥}�\#�w:ƞD&�ȧ�@��M�xF"�1��*�Ԋ@�蘅�8ꃺP"$1�D��A챦��d�� �0��S��GO�D�� `�_�g���0�~R���5D���D�!�1=�1)�N#�
�E�Nk�'xʳ�J�D�Mn^!�W|��S�P��ɲyVU���/�R�{���~�,�3(y�m���g�)�|��"�^��v̟�c�J�����һҖ�����s��؁����i���2��@���'F����;��V��j�l��}ѵ IԦ���nMsοX���9�8�wp \�=�FZ׸��Ȏrw����%֤�h�m�A��N���WVo�K;�}�����9T|��̬}F�{1�4!QHՂqH~v'���
P!�N�ޠY��Տ7��d�s�U����VQ���mgGS~���j��p*V���~i7��=a�f�	�4�M�f��X�:߮�nI�H/���|��_�߻k�[{0�$�F:k~���^~�@zק�r�zN���2ly��A'�<�f�����Ĵ��;C�
��R煎�y��equ>ː)\~�=9b��B<�)zѲub�o���.l���4�9��r�V��?�W���%� @�����
SRU�\w�"�Eź�嗴)�S�;���n��׸�_����{��\z��<Q��@�Ǐg���H��O�Yv|����4��z�MN>o�����B���f�k�wbQ�v+�g+�P��4��؇�w�V�]A��M J698��AZ�w^i���i�G���n��?�?n�Jtl�
��jXa�cd-�~�йzo�[tbU!6H����oG�g��, *?�'l����r��
lZ-��0��k;"�S_�m��7	�]6U�p���Y:�C�Z`̂�Y���dM�{�f�
���N|�]k�ϧ��"N�ju�^��z�	�ް}�������-���qV�V��}�o�z��K��Lݸ�e$l��{�h\Ț�Fj2����&!7���赛g�����x��*nc�����DƢ��"o���aN&*zB�!�V[gA��é�~��&�m�]KձA2ۓJw
Q�������O_6�/�&�~L�VB�Ť�XP�n�ѹ<X�ud1�Ы烶P�W�5���ȃ\�%[h����&�i��Z�.�V)����/8�w����l�Ǚ�I~�J�-�d����*��":�/��k��pA�YN�C�Ӡv���l���8��oN;g�i�v�zy6,p��K�8.�a�p 4�4K��S=�J�����>߳&SM��ݰ�*�O;5I�j,�3*Θwy|���?�4��.��/0��m�r~�o�;�y|v�~��> ��= �ٔ�Ïe���|��wG�S�u����(�B���ς�ywV<��E�,韁e�~U��5��w��6 LR]��T�yf�%C��H�HG�e��D}�T�H�Lk��u�x ���!&����#��4�#?���sf�d�cuA$z�	�S$�ŭ�(�3�Z��UKez��-�"TB���P��,�����8���AΓǀQ�.�s�����1o#������I T9$���=0�:�R����]L;>��F�)�F|��em5,t��~6���G�2LY���y(]u�C��C6ʗy��g�3�:�36��cԏUm�Yd�{��.���e����I��݁dv���vc#�9/��q�|j����nQ���Nht�Qm�C/�SA�R�*�{�.��Z51%��y���๓;
n4�-�oE%ס���8<U&�ѵ X����v�:��?�ol|i�M����o5�-�Xi�{�LT�̚Ȑ1c���Qn������'����^ f����o�`�_ߐ��[@S�oas�2���,I������s��X;�^
u�٫F+�O�Z5����*��Uך��n6��_��$ ����a���;h�<�@�e }�7w�vF�(&�W�'n��� !��8�jp�����A�4�vˣ�S%u�����a�tFwX���3d@TR� �eT<��|�0�O�_�~7��b���S7x!F(6BÖwB�מX�G���,�b�,�B��@��)-��ه�z-?�JvF	;f<����'e�0�1YOS5ak5px��x�x�8%� &�lV��x<��ۅ�C�"�/z'H�`��^"􋑬�F�ˇ�,�+~&��ywc��x0�1���|���'s.6]tf���^�܃�����4��B�q��S�W�2tZ�3��ߡ�-)��<��ιqB�l8��/gƗy���o6@��G<�d�Н<�Ot����_��{އ�oPqP���AL���	�Dk٬+هA��C��"��5��)��Jj�m=\�D���w�8��Ė�ߝ�0eDo���P�_�H����Y�n aqJd��J�6օ�~��(���S��fԤ����Χ�($�P���^wb_�̦���I9�ǹ�7����`;h��%�^�$���z��������۞�٠!`'#�.(|f:���ʫ�������PmN����]8n�݋y4��W��j�4�����O�2V��*�v���\af���(Ȓ�����:n�jm
��
%"�b*K�� y�S����Պ�y��|��OԞ�(ۓ�H��k��[�`�/ JH���s�A�C��a�*�jX����_��q�6���QJ|_;_:���va9t�^����u��,�E_8(����P�.�l�-զ�pf&��r�����ԓ��ŷ�)�
z_�A:�@�l�����/��~x��+�|�Pª|�'�xg��h��������|��-��RD�m8��0�Y2T������~+s��i��u�>*��z�ͬN�ZJ �򈠔h�\�Y�5x$_�ַ��o}3ч�8�?��\��+M��ϷwFB�v���M�V�����1���T���F����U�Xp��[�O�tU�+�o5�as}i��1��� B�o�J(��O��+�²F!ҳ��A��'��5�}G,:�#�K7��1����ﶔY�#�< �$�F�0ZS��!Vv�ȔB�8kx,_*���Een�G��N��h�e��4�!�J���D>WU�>��fSw��4���V�3hF�]�����Hz��~8�?R���C���)�j�
(⭉��]��$��?��B��qM�f�g�h���ެ�8�T���D+�fߝ����j�K&�c[9�Y��S���s��1��� T��>N( ��'�$'��z��b['����I��'���Ex%؉o8^U���ܹ�/�?xCÄl,��k��a��O�C����j!0�
P��O�n��[E��Q	����O^p�䊖'��y]�z�"�����o2ơH�c�����Xq���b���(e�b�=��,:+[s�L��(��s��S�g�0?K;m�[�EUV�?(B��I,�<����A��{��i�i�!�,��5�y�|ߵ�a�~��~C�hd�F`�����'�ku�r��S]�2�;��'�!���ֽ�m�ȓ�#jU�ֽ"�PΔ�}��'ģ�T.�8�^UAX/�ޙѷ��b[+;]u�sx����2��~���48j�>�Ebc�!�#�>���bUiW��몑4i�����⸲%�G]���Vo!��΁��R���D,c
�sϽ~�%Ȍ{�k����?�T%?���Q���:�$A.���}R�)���lD�b�8l����G�|qR��ߛ�ވ���y��9_�0 }k�)�+*�v��ÈY�@E��N�K�"�	�tR�&�Y�^�۠|rD$J��|��H�퀌ɿ�_����Q���w�l;��7>whS�-H�Q�E��eۗ>�!�m��N�&ↄ7��[䐛�&�=ah�6-�|M�[�E!��>"<��|R�Fb 7�,��$G �u�V�<_,����P7���8FZ�P�������;�G��	. �F)!�̮��ݯW	��4�G@M���C ����ѠGO��":��6�ߒN�@� h�4n*1�m�S�=�gd�z��I��B\�,�E�|tW���7�_��q�'�cA�.���3u�QF!t�g��Ex�ג��3�S�e��6^�O��
?o1V��G���7�䁂,T$�i}���TR����F�g]I,[}�����Q�;�o|(Q�.�Y�O�:��E��sWS�G�B�Y�R�4�B
[���lXxIr�KI>膯��tc\�f��
Ë�$�*��2%K�e3��a1L��8<��'�NM�L�����i��§�|��a�ϤÂ	ɪ�1���>f�Z�|�~����-�E��G���+4��I,�,����a��'~a~�e��x`�/uk|�Ǳ�&-���~� ��P�!YL�p=q��}S�����f��ߢԌ>2��Q��� )��P+�A!���1���U��,�!��{��'�۪�����Dn�)�m�5�������9��Aa�:��b��gg�I����҂~�~�������-&�����.-�Ƴ��9@sZ�4H�r^�N����Zzox������U�#y��g�Dcؔ��¾ƔH�;��ZQd��y�A�����P��T�)��L9�s�K�x�+V�Ա��^�>^4��12{x�Ws!x��#���Da���L ^�R��(�� ��&�q�A��
܌�'.<��A����zk�22 �#q�3,�6u{fJ�ݒs*
�2V�Q���fh���ZVe��(�6�Ӕ�j��]%����C�5D�4=�_�+A�]3v�U�<��a���H��1�u����%&|l�2�-�~��Ώ��pWjz���_Ƚ��4*B��Ծ���!~��D��o�������$�F�eXZ�����Aa���E�� o�|F6�/�吋yD�El��S#�{����IV���+������y$�yC��77�M�Qkw��X�(�Ɨ�Оk���	2���U�%G�4/�#h������C#ⷽ'�"�7�GΘ�~Nz�a�V T�_w{���C6�ANS�-����vi���Xέ%?L���_g��M&��[�]�`�%ro|�q+$вJ��Y�1R��@}�T�����Mg�#F��:}�O�R%N!6�����[������( ������o5Ʈ{M< �`5�ɍ5A��1K%��ȀL�ǨY�F�;��0��R�341�g�Ԭ���<��p^��v�8~���a'��yyҶq�ʎ5��2 �s_}�U����@��;KyK-��圐��h���({��9Ǎ�ؑ��)��v�'���ڹ�rDF7�P���n�c�öT6���͵TX�}]OnF�:��Y�ڥ�bl38�.g>^�D�䷁���6��`"h�&�˓�C�XT��>%q�4
��	�6;�I5��!2c��哥L��R�eg�(�#C\h���4�i���k�oY�Z�I����+s���u���<P<�!h#��[����U����X��r�|KUV�%j?
;bz����*4~˕r�y'��X�W�q��h5m�ԩh�>n��R��CZ�{iw�LiP��	z�Y�������\�@d&�7�>1gGee���#���~<|�ZR�B+#*����S��cJ�D�GL�ʯ��/UCe��#�i�G�����i��GG/�F��-����g��X�������t��k��=��]"�������@�c�+���L��O���x/g�3�
�X\�� �F�4���	��Gt���*�R��eN*������r���2rL�ω��J�����C/��z�"݁S����Ja�M���2U�z�R���;k4��hOXW=Z���=\!|�˧�%��6՜b�/M�˰�j��y,3�Fh�ʉg��5p(M�Y�:��Q�R�q�H�ѕ�c��-����A?���$��
3���ɗpL��P��'w_y�N�����%��7��R�R�}�����T,��(���MVu d���ѻ���r�`�{&� ��G��z��r)Y2[N(T����^��ӹS�0i��M��cV�7��?�Wg꒐�fRAO�ኣ���"F���E9~2)4%��U��4u+J/0>�{�S{��eI��N���|,��;[,�&(Ȉ�;�5{h�@]��PR��2l�)�f��	�£^��8g�^R��e�2ԭ�r7�����8��[ ɪ��{�3�$�f���ɥ|#�\�Y���K�ۧ�Y���h��U͑#]芇_�Ҩ����kֽMk(�ӁeJ���D��n�]U	�ƨ�C�W�
�NvF�z�c���?�J$�����uhp|�:��xYf�Pܜ�N�;5��;��@Ҹ��1�T����c�qb�p�ۥ��_* ����NW�?�,��%��~�<�
c�����=�H]�ݘ�奈���6��s��e�*k�Q(�Y��H;�U�>'��9u����ˍ�Y/�{A"J�x��{ЀY�)l~���f�Gs�Z�8���4�*�x�$��AHk�w(�F��(�;�	�,d���J�MI�^Ǳ�E�"�?��v9��l�PʏM ��㻽�Y9i�u58�1�����hxDa�)���z��w�s)}���3�>�&���8��Ŧ2[�2�U���@,L����@L'쐚j����a��m.<lG����a=U��u��{���N�O�+BB9��b�@��
�{����<�b��pp���<}�Җͬh�á��K,�?��Ծe��1̗\\HiKA%�\u��Pe̡eb�7҃'F�� �����B��Ԍ ���US����Kp|R�R��hw,�Bp���ņ��4l��;��iG��^�,�V�8�5@e��G�q�'����˅x�Ȣ��t)Ϥ"�YE��R�.]�B�����°��S\)��Jb8 }�*p1䦶L������k(1c��Ƞi��V�ܖ��f��(�ۭ���ԕ�r�����@�_J�'�3bwv�Ap.�"����@�4�	��躐���ؚ����N��p<����
�p��jU\�������iX� 3�ψT���]l�,�	�r$�3/;`�S�1��t�֏CK���L��Pԛa����<&1�]O��<.*rԪ�`K9�%����t���Y#��SݜIZ)`����@��l�!��ĽL�F��Ȅ�W�.��"��׬�)�+�iұ�1$U���>16K�gAw� '\��,��,^:��C�U���ց܃�U��QV��� ���=κ�A"uy�/�U0���m(IPF�"ݪ� �E�+տ�Vulr���=�s�!Ͳ���}	R�xa��
~�P�d��>i�ŵ�a�H�p�}
zۏ��z2�^�p�	��⋣h��2D�t���x��_���,��j��i	� �?�e�dN�a."�� M���*����I��.��l���F�L����iH�]x��{H��ld۫�T�֔<z�ʜ���x����^<	
3�0-Di,����i
�ǏX:\%u�E��*��,z&���$�9�}���{*1ާ���6åBRMGC�Ę�a��-,���[��i=wh��x�Q��Y\
h;������ ���!u�������3�B԰�u�� �-I/���hL��;�ۆ�-=��e�qb����$�e	uEA�i�[(�B���]��,ćo�6H��!,*m4���+��|֍���2�P��Rw-(���Ow�g��NǛ���jRю��������7޸�h>J�h��F+����H/���N}ıv��S1-	amA��,)�2��j�L h�h����9�Kz�oЋ�3n���5`O��0\��W2�>�Nj�/��/���DWBI�Z�R�J'���A��`��rhԒ%Y�)�Ͽ�;������3E��O8�x��Kx>eZá}Z�Pr��Ь����S�5"���$�Yw�'A@kF~Aׯ�,ʬ8�H���<I����O��yC��o&�������
����C�߿mSM
 4Y煃
���Fp#V��'M�"^��?�����~�PE�*7��LS��+��+��j��\��m��:[�ٌdj�`��;b��t��7X'�w!\��s���Ar���/�� ��UtQ�a~^��SR0i+��Ƭr�n�=���YPx���&��Z��㦻��$3�`%����n�}�Q���/ETb,����:�j�jg��=^��w���.[%Nٙ߮�Y@OV�Opr鬆)'���G?B���fP˰��"��Q%˲`٥S#��?�J�Xr}�E��Y�'���ۂ+jǐgp+��i��O�ȩ�s���\�3����<k˽�#��Z�����?]u���6p�|�07�+8�ƅ��@�@r�^MoI�m���K��u�l W>��	Eh�9h,�����g�b<-w�ñ��x;o��|�Hf�Cn�ۛ�Q����K�@�2�cMMƬjrk����s�M�,��∥
�퐤�I�f����r-�"����e��B��M!���D�a�-r���֐�D$]�IPd	�tL[k�?�P7{�	����#`E,l��쎦�$��kZ�bI�6���i|�M]�t�7��g-{�-���R�ԘٞP|�Jm;� �4�v��`^��;�>L��z>���7������s�YKo�k�Cy/�:D��\hY'��(@�x�t���Hg:�<+'aoC	3�e��169$��p��V�5c))M7�%D��a[S�D71�x�lY9���Iw�*��[2$��$���\AV���]��H��	�l��߆sZ��i��bϩpb�I��Z߅�
,e�r�o��qфh�4,Ud08�L���L�R��"w;���9� ^�;r%�D���N�S+�o��V�Y��M٤�V�y��9g,A�cڙ�`B��^�kRl�����e��	y&���Rp�$�s-��Z\Q9�"�:n�K�7.�ݰ솏 {�Y+>���wa�����\}'/�|'�H�Z�$���Br�E�x�\[��
��{c,χѐV]:&��rQ���[��}�5/�"$�Ē^/S
y�殎h�=}��ɱ�v=�7�]7n��H�{���1�В�!V�U+��v#tZM�5�@���D8�?D���7�[G���\�:�ī ��(�H��M
�&Œ��h��K2�WS��1Y�+&��ŵOgI�QL��x����<EFc֪Nz�	��
��h82�L&�l��õ�u�_����j���/�[dbuV$�?�eWC�~Z�1<2�8D�F�W�q���	��#�B�
�rgIb�5B��yz�iC����?!�~�(�y�kz��<>��IO���o���Zغ� V��h�}t�u����N`v{�;�.+w��S�4.�aV��+@�w¢Z�#(҆}q�mf�7Y����������b'ꔥ��]۾�*z�9r]���UѝpS���F�5�(!n��p1�Aʈ�eE�Wǟ�
����
i�X�j]�e�n�����J��v��a��U��x� 	��Nq$?w��0�ipŹAݐʸ���wg������kWX�~
?�#�����P7�;XW��~��:��u�Jtl-�)DaӁ�y�\�kc�?a��̋~�����5+��K㹐�`wy��S�҂�@36����i��`oǏL�c�CT�]ެx�Ǡ�fJ1�I>���:H_��4�����u��q��%�\�h��rL�D�
��RG����� =�<��ڧ0��Y�"	�?�V�I�ң3���3�(�E�$/�F��H���vh��pmZ�3���FXA��`�<�p��~�F.��A6��10���������#N>�'K�9��Z�Rچ�;#�H�/�a�0et����u����P�C� hN���q[,�%\�&�ıYh�����W�'��h*�R>�*��˽��'��*��Xc�!���Um��$(�P2R�R&P�|S�G�n��ƪ�1�����[� ��e�4���-�8�kD$H}��{�²��td]��_�^��hr��m��-�'��?��<�LA��ۚ���h�b��wL=?��;�I�l��F�pE����ظ���=�W����B$(#YX�NM��v��+1�s�Q�buzqe�ƽI=��([ ��ժ���C.�H��lu�6G����3K�:b��uȿLͿt'r?yx�W���QYР��α���6��g��%�@�lm��EҺ����C�m�b�vG�wuq 5��o0[-#��V,v��c�@X���PTcJm�l2���Ghk����Q��o7*��N����2^4w���#i�xn��|2kDl�CCŊu�A*��1�����ټA22�&��-�~���AIx�2:�?����&�'�QJ,K}D�&��
�Z�qEE��`V׾b�h)Ӵ�� ;&�We d�9��r��=44�rjd>}�\��8�萏��s�!��\��+wZ:�"��,-�媂MUI.S�0(�G]�b)��1�C&�biI��s-���*�ά�H�n;�71�����/}^r��ʾl3Г�e�u���r�>������Mrܸ
e��Jo��k*���fV��*"y��Z='M�:�K�;�ۤ�@.��|�jd��$�F��N{����������qĖ��{�d~�t��+88����} �ش�G���\��@��^S�a2���<7ee�M���ۓ�L2��O�Lt�%+��(L�m
T�ܺJ������N��Z�O��C��%�O��],Y�?�ηهLV"�=h�-vc��6%�&��A���D��`�{g�s�ȍ<��N���C����ĻKa $Sq��mvM���ux��Q�� T��
.���ဣ�D�,���@����]l7�w���5p��n5M�c�yrn����]c�<�?���chK��[�%�{�T	B��xv�	,�����N�j�Dr5�Τ�geţ�v�$!±p��j����)�؞��V@�$)��5��̊h����~u��GPk:LEҬ�Fv���!B�oEހ�'][� B8\V�nk������������_Ҍ������^�/-���w�8��2�7�qhnwUuϲ�Q�u65���v����ۅف\�ɨ�� ���-�Ğ}�ZCOx���羗�FX�Ґ�3$ܥM>cN�����Ę�x明�՟%��º�\�u�M��ݜ��8[av:B�c��vB��/�~ρ`Qf���|��q��V���DoW,!�z��΍`v�t�4m����l����/��G�W������,�S	�!��hJ���o�̌ݾ�ZJ��N��k3}��l*0���fU֘��I�����@����H[b�P���ʔ�!���q��2�`�txp
To&jT��R�關��J�#,��l��R��W�g�����o�z�O&k�����E���:l��2S-�̽ֻ�0L���0��o���-.� �MOn���[���3�b��(����0 ���Q�!������l���b�7?d]!O�%�3� ���e�i���Fu�)/L�RE>����Z���u"�La���S����4���dtZ*)nz�$V��� ��X����M.�Sl�t	[�r�ʺ�8;�rȊ�ƭHZ89�ug�5*�>��|d�ܳ�"zī{���%�ƶO�EJ�q5��%jA���٭,!�/�k&D��0U�\Z(�Bͽ�[\�*�L�ZB{�[�(�K�v����w���F���(��A��%�r��Z���M���%4�Bʍy��o���:[V�^w�f�£8e�3�� ��I/������,�P(q� ���.qB�9W+��Y���a�V�Ԋ�'&x��,f��J�uX�V�h�ѫSTk��b!h	���p��tĺ��x�#�U�cR�T9rJy�l�b:4��b8=�4'�η����a]�K�)�9�b�Ŋ�bh����?�tVE�[�-���Wd=_OZ�k�{"qv]KJ%&�����!�+�Gd��{�۫Re�{���ݬ�4}�����L`pN� ~�hw}*T��h�?V?���\�o�ڃOl~H_�@��0:����D�Zd�"�v��*
����>�v���XL�W6�~k�*ޝ@})���Hjy�-��`�G�χ?�}���t��U"�{���,��q��P���N����F��� s����7�j6uY4�������=Ȁ��Tڂ�%hy�kRC�ȱd(ަ��.Xc�������1D�Ne�̐�v��|@��v�}Ee�&sp����æ���7/�~������=nU���h����wT��]�L�k��u�E����Xa��#��xb��ZJ�j�(��N��e��~��X	AIb�ޭP��+&�L�v���m��\8C�Y�Z 7��B1y����o����
�6]�ǖ��C���1\;IT��u� W(!�Fi{2w��h�`�V.���n��:u9�I#�}��3U>vP
z��)͛�ҙFM���,w�~.�8����oI����c�ؿ����0��S?�l�N�Ӄ���u~�2!4u�ƼvM��Bf��ҟ'�̡��p,��l�S�k����[��0OY��D��3w�<]6~ۉ�p�d�$ʸ����O�Q���͋l�,�u����*r��c�$�U}�)D�\���3_��n{^�Y+6�6�ɸ%�;3�wX�(D�Мa��ѠܞTr�=1\�Vva�x�NQD6���ruӹ|o*=�e����n��.X�U5)�H�ع��KY�7O ��(7M#��/�x�E���f��&|�h�G-sM�X��.��0�wٞ1���@�/��03j�!x2S�$R��E�OO���lE1*e����U&�	A���r���sю�8�}*��j� �
��tr�d�gҙS(�T��8�}��W���Z�a�6�F{-��6h��^�F���4����A���ӡ6)o͞G�Jk2�%�pҔN_M�Kճ�4� 4'�sʑD�e�����>��s9��ߦM�K"�S<wF՘3[��|��]�_��p��^h~�	s��.�ҷ��v�A({Ă�<֏zm !>�k����-"73�~�D��wk�@u,�7�X)�(���gb�!�NڨE����_4
�{c�|w Fo��b��E�,�:����b������`�|�F��X�q/��T��bu�`VM�eY�\�{huF�0�XxX�P�[��8uDa\:�Z�����Y��Z���u���rv��t�/OK��b��$l(gI�<.�C)SJ�rS�q��j�2�����`�����7[H����jp{�q=���b)}m�aD�>�r���cc�j��K��7!�������aMo��j����:���/�a�_%]�V�:��/����yb!9�悈k�:ڢ�̏�řE��~n��TP���	IX�6G���RyY�W@��^5A��Q�2�ȡ�ћ���|�&���Ɗ��%��LJ0�W��i�:�o+�+��d�_�S�5U9����1���#��QK����~�!km�ʒ��� FԳ��<��̎�Q�N?�D�BJ$sy�`�B�#��8�A4x��sb�|�n�L-��(ċ;6+flA���Z����J M�ZKH%&l�uh��3�$'��s�� 7����P~KQ3��y�|�P�5��T��^���`���v�krtp>��m���*�w#�6�Ƃ91���c�Q�=FU�����[Ǿ���p�i���f�ym�U�c���=��CZHF�l�f��t�
Ȁ���Y���K5����0�,���#�e�8��aXg�h�4RFqȢa��вA63>��Ĵ$H�F{;S�笧�Z ]���x��b���M�t5KvkqYc��E}n�2���H���B�s�T�F[e�Hj�T�L"�?ڜ�+;�W������W���ͼͶ_��mQ��Yk��8��)����QMi?�v��|kd��9����-��,{@����. .�-��V��X	S0�	��dI�kG�G��S1��k;�XǶ����_b��xU���C��/J�c!_��-굚��$9��	!���8���'��c݁O����Mb��/~=�!������������������x�1�A�PI����	���<z�ۼ$�X���ʮ�)q��n1F�(�'���v�k����c�Txu��퓪NUv�}��@�t���b���H�$KDJw��P����ZA&���<�7�0����0���*� ���-�})>�j-��_"���KJ��� �,7���_�CeZ�����9�HAn�G}�6	�̂q��K�M�@vO�H���C���Mp7��z�9��-��a�p}�H��0�巀���6n7�k2�X�"g�.܆ 2�{r��XT��Rt�4
��m�y G%�l���ɉ����D�vtU�A>��֑$s�ӷ�t�.���b��]E��`��t�@��k��Q�l&��vv��f��l��>yy+��L{U-%�W4 �i%�=�a���E3�#�	�$��s+�\��U#~��+>�_)�����E��L����Ӻ�[�6hu��Jo~��ݴl&�ݖ�&rp�x������D�s� ������uύoꁭ�<K�y?:���fk������b��b7�;ب�X�E6�¾C��ݸN�k��V�\�`I-ʑd��]D�d���5g�tBc̿���
TD\:)��`�Ƽ�|��A�[��]/	k�����.�8x����&m�h ,�P=�~���WBg�5���y�����3C������ڧ��_��s����4g,&%a����!W���oM�p�<[n����a�Ib�%<�s#)�\�f�Ċ�2غ��^�?P���!0+qu�L���T�����/���oU ��P�V_��S���sW-
X�u�(͏M~� ,k0�Ak�z�T^@"xH���G r�}�:���n�01�H�L��:���!7��(�|�b����mm��.���
p��QQ��I�*��2�~�\�����[�Yjí�����$�ǝ�E�󞢑.�j�s�4��"�Z;�	���w|��)1쏱9��M��N�g�Mt/�f�j׸ѦS�G�V,7����Hl�Um 3b��A����{C>Rw)�6�+�I�[1��z�]*1%�� C�:�\�m��n�w��<��'��Y�C)�!U��(�ª��,�ב�G�.R�"��F��}�ZX��&{�/oˬ��֮0��T�HK�Oi ��"e1mv�1ʭ�!p.�ڷ}>=6?Jℒ�п�����/ĕ����ξ����Wa4z�O�����W�����r����&����>���G�A��5��Ǉ����ǎX�)b�Ba5���M��v�o�.Q����..,��i��-C�3A�2�^�+"�4�Z���_���v�����l>[8�;�B1���\��bÛ�.B�.Sǃ�*�����i{��j:X��B�X�Phd ����KR�����&�Y\`;�|
tw�¢�7@e#��zIԆ-+auV��!(��1���s��ٽ�ā����[a�z_S��^�䶘ņ$��rc�B�2ހ�i�_
N˃�Y.y?��Y3��4Tk#?�@h`,��ܹ_���ɘ,%͏(��;��������x���Sq���;��-�~<���g�6��9��!��qqt�VZ�Q�NX�c�䖦8�̡I����.����yh���u"W$�՘;�C�@\��s�g\{��,�k�}��7;��gZ�� ����G����,�e���S�kp��%�C%���(?�V��zM���^���S�D�����6dkt�>W�D�
mQ��E/P�p��5���\�7�������x@���;'����@�;&**c_�
�\���2��g�cD
]K�6P��kSx�k5ԧ|;�l��W�P�r��C�r�fJ��3F���{����3�d���H�/���� �#��+c��5&�����c�v��f�pk�2S���Z�I�Ф��-����%�/��#H&���{��>/�F��K��{\P�Cr�b��/�9����^d�a�R�;�$s;i�k�>8Be%��@lf1aFŇ��V�;�XҦ�ߘuUY��yƬ�ɫ�IV7ѥ�.��`�!`Ri���0w�ͅ��:��x������_��&�u�L3�B8�G��]m,+�Ɂ��QTY$���0��ޜ�Yi�GG%WA
��O5�g�;�s�cۧ�"n��3��m�z����Y���%йLԉ�Hy~N���H��sZ��{�s/�/<�B5��e2/�K�%h{I�oؖ(��BMuj�yx�EI��]?��ڐ��K`ag/�C��*;ٕ��:�v��r5K��F�}�l�1��F�ӿ=�.����#pg�\,ޘ�)�s/���v��¿��yR��L��$ъS�ݵ`{nvױwb# �B���
a�Q��Ą��X�a��Ō��>�4����j�B4�-�����|�Re7�_k��6�qb�م�oh���Y�� ��:��E��^����njЬ���~�N�Jڀ'{	�5���ae��f�h�Ǽ ��R��pB�&dT}Z���=n��{J����F�]��o	�m��^�v�P0
�0��Ȍ?y�#"KE�y�3����@�]���`<��x�閷,��m�z��'c�b�E��.����e!��2p��V�!ը�JBď�?Pҵ���U'$E��b�
��^�y����[qpF������!%3�ep��q9�{�g��H)��-6*Z�L/����h���2a�0k�k��v�#;!`�����4w�P�mx2AKI��n���9 +�2��ƀ�s��?�>� �\��/��>��h���]�o��RK�=����M:�����ҜR�����4",4a�i����bS�}�6�!�>J�Zgק�}��'�|�Dp�G���4#hܞ�/�����Q֌����&�J�:�X�4���fSSq6F)j��B+A}R?�+�&�)��[
vi��������͎G����M4�_�97rcW��5㎭Bm�:���B��P %�8+Y�+>&�E� '���g�7������SȚ��.�7��2RW�XÏK7Mv�k4F����gA�sA>�(���y���DOF��!;���]EjGS��l"��i{Q�k�X�������pZ�+	��ʑ���%�~�Z�㱑� �%��[]x� Qߤt�� �͠�~a�� h�AD$���9/��x-;�N����SM���X�sO�D�_�ɿVJ�>$�be��;;�%��������}c`y���'-H�>&z�v�z������ӂ���#�݇r3b۲���4�ŝ��_r�9�hgv��a�,�>��x�D$*w���(�8��=fP��U��8?�t�V�g�퓆/+��Ԇ9�Qݣ�`����$e�+&�iԄJ�:y��S��͉�H���k��Lկ]�SNN�eO�G�e���W���(핂���i�=�W'�>�vex�m?x���3�;"Cϰ���{��{��=0C���W�+�T�}���������B�u���9��搓!,��F?�����zw�l|��6W}7Q�z��Wx�B\o�|Mr�q�;���?vI'�`���ڢ"�����Q��K*za�< ���������k>m����9ihu�1؉������l�fF`5CÎ�2�e)M�i�p���v��E<�v�19V��\�NQ٨B8O�M���6ɵ_.�؟���[$��s�h��!�n0�l=Ք� j�@D�#¾�f��wZqϹVx;�⬟l!>u��gs����q-#���[¢�`�IN��p��
�d�F\�z�c�0R�؏{�2Qy ��S��
��
�\�'"X\fuV�Cr�If���_=<����p!:�	���/�"��jg�:�� ?�Lؠ�F���,��a�gς�ߊr<_'⫧���E�$&�H��G��֯ s���a�̙i=�g!a���j��ƆDx������]�����	{����Kc���ß9��!���{�j�V���`�V4�=��B�I��R^<,���N��!���?[��o2�yC�Mr~s�>$��ec�I��;�-[��8��'�H�ڠ�0l:u+\���D�M�}���uY�N��������o�㓷��IQÔG��o���U�Ĺ���e�;C�DҸ��`5%�}~��գ�G+ȇ�k�[�G���	�y��D�*�p�����bp�,���m+��+Vj��2M�"��<��;�fRl�t-˃1O�e���a?�OɜU
���N�^<4U+eC�~�!��t����.�ծ��x4�	��md���N�ҹ�H^� �qvA�,��ִ����`M�2/�
ԫ,��l2���x��/Sk�h?K3�����v� k�]Pu������׃�+�Ov�_��j��X�~�M�ƶ���-��*�q#0��R���G�?�������9MEh���NhsdA�}�.)�����,�]ȋ�ں�H>i3�"�Θ�ᦧj�_� �Z9�N�����j�,[땵�3x����<�N!ϳ.�L^��GOB�Ɯ���	��}�
$9��\f({�	�#���]K:ʟ��*���AY�X�c�ApT)�ٌ��-�@T���=
,����ɠ��%��SL֌ũr��Q�����a$2����(<�g�d��X�>��/��`�iA��lN�+�<�sGs�Z�4��g��z̘
�:�e�`���.��"���?���>J�./'v+�t�w�y�l"�G���]�����	/�ש��a@.U�@H�I9�� ��>��4�2�s���C����\�X�M,b�}Un�5~����-�x#W�׫1�c�������ȩJ��(�٥��1/%�ʙ	y�U�R�I�Y�*��e������ѫ�`]�-��M�"V�]�ށ�'�g^�@:m)T���9,S��O�yx���J�E��;�07�'$��,�I}{[B���0�>�zu���Ղ�e>+�l�n 5rWX��,B�A:�5�������l޲g�H�������.�!k�9Z��[kו��w?oN%P�[/m̳�q�X�;�����������3t�^����*�<�\p7ov0������6����z�&3J���z�!8�}.��>�Yơbd^�ۀ�βh���+łK��E!80M�p�8�!��m$I��.mh�Hp6�e���P�t#W��^�>�g�[.�^�����n�3����o9�͠bE!����#J=Sx033�E�%V�|�K�+qa3S���=�JM<��;*n�b/?.S�)�I�(�����-�����Ͳ���	�󷜻N�F�B�w/蠦e�<f��������������$�"b��6ě܊�n���t�I�G[�b�Le���F!
̴lPǗ�yT�El��V��ZzF�3���ķʲ��\D��j�������i�R\D;�i��3/��p��[u���şne0�k�V������BG�$eӶY`U��\��,�/����w�O���6��B��m�kt��7q"����(�&��@������n)9!��Fh����"��eI���n{��\�������^8�������]l�&��U`���vSU��}�/I�~K��S�F3L��9b�Iڵ��}8�J�O����B�\�h�9����42��6��L,2w�K�\���M��RO q����r�Z�+�Ai�4���i��F���L�~��.0ؽE����Obo�6��ɫ�̻�	���)�`Ȯ�ؘjhr��X��{�t\IM}�0��[sلU,*m}�v�����Y9�yGYi��0��=Dvy"�vX�^�^�<�`���� Eמ����(�����V�PR`��\� ����F�Yw��E�fe9 ��u��xe:�)����B/��g��8����@�	f֮=R���߹;��1$�5�F�N�WWK��4���Z^�Sy�F|�I�[�P4��O����o��[��5O�`�����T9	��04�����8o�q�ߐ�&9?F+ǰua�O�F;��uފ9ux9@��1&Lx��X,{�p�~Ռo�d���`�Bd�C������O�Ț��ǯ�3�9wF�2"axƻ �;���.yzփ�"��Q���DB�n˩I�x�� d~�N8�/�1�����ḷ�4��|��Yr����@o���a�#9��_�«˖'�3p� �I%Mwk�@�5�A�\��ޯ��Fê���?a����J?�)P��>�EY�πu^eK�<+3���c��g�>v�^H����x�֋���c���Vt���c�FU.(F���|�ޞv��0�!T����^�&&����D^3�D�aK{Q�`#+E����b�i5;wx~,�RZ�ҳf��8DH��l_�:���,�g�(�
���� �g���9Ԉ�ޗ��	'��(�¯�j��P@z�h�� `�	�}N�:^�0�},j\!���~�u�L�^2�d4Tz(	��]�r��j����Zͦ�Ҵ��A���͗i�z�zt|�V� �E���4�����\a��!�W�t�G��u���ah��῎0C7I�K�I�����5k3�e��^�f�^d�[I�7Q�gLY�u����嗢�j��pC����ڿ?��Xw9<5��d���?�¿hǝ����	��J����%�yj��4 ���i͵m1�n�1�����>�ݿ�!���a�?�v���t��QcW���������Յr��DlT�8�9`�����v�����.�dp]e/�a�
����|���qP�W50q��G~{qvY� |��&��Y<�9ޣ��t�1��ol�Xȴ���ռU����5Tu��薮)��@������ZQ1E��{�9Q�����L[�n�T��I#B�Q)u�Z��u�H�x����=�����gj��g��{����DD���$e��ÓЉ�" B8 5Ǥ��.�lJ��v������DS��U>�5�z�Pڪ�Z0?:�=7.���6ړp�MW3r�E�N�E6t�8���^�dX�Y�1ێ�����4�B�xJ7�.��0��,&a�����M��9�&�t�z"���t|�0��*��|D��=�d�n�V瘊8Uf`�OU�����体�:a5���_���j��#��kQ��A�{B}��0���51N��vl$�r�-�,��Y�v���!�۵-9���̺㰚�U{�f_�]]�'oWv�zRd����{A��2Y�vOm�I���E��������hv �ier������e4��`���9��p����W���f�P	����,�v���~���7ʢ�>��d�Nٛ��f�x3]\ ���P�X���(�F�$c�y,[���Ԍ��gH�;�/�Gd�Gh����tj����!��y�b�JGE��q؂.�R�F�5���p���c�E'�<qct��Q�~�=P�O�3�� ��d ���9Qwo��i����~N����~&���de�bD{�+&dD�;�uV�},{M7,�)��=|D��S�>vT�r�V��xd|�[����Z�0i���LTZ8˦!�E�2��ʰ��'\�T-*���:��̧;?���=d��;\3D �zb��b����TX_0���4�OH#�d�m�&1YKD���ت. RRd�$�	��V��S��>���΢�o�~O�=����*�4o]Y7�M1��d��O�3��}���Tr���`�YB�!��? Ks��.�LS���^�)�3��q2R�踱��[_c���Sr�^ג[}�j�v,.��<�Yҵ� ��ϵ�=�@r�'�� �j#  �[�)>u嘩�Sb�L4XR���R�w��v�����y�a��%�4I���b�b�N� ��8B��oP�8�;]�H�=Ah~s���cF	u�evtެ@�h�[��H�Ig�bx%�myx�9 "��|0�u�P&H$r&[�e"~7����i/.ï�&0���xU�H�"]z
She �*�&��5�R�.�e�x����D%���ki�Y��TChh���-��B�Aw� ���^aS��%�:�mj�1�
F�&*x��Č�2�}f�X���MD�Y��0*��V��L��
��UT稛�����sļ�s<2�m�Xfy�,E�p�� �"��%&(��;#|� ��
yA{o���W���ZV�a���,9��K��p >6lj��Ue��iZ��&J�ଇ��#�&Q2��H���c�%@7��V�>]̓���y���@`뵑�����t	��WD����c�i���.����-�_��2d�9}M��ƴ�+���y�q��4>���`�?NZ ��÷�:��P�Z#ZA|.�m$fӮ 	ܯ�D.�vc&I��}�k�y��Y+����SN�7����ui����Ƣ�$a�
�N��B�\�-�V�1ř�6g>��Y@M;Z�ɞK��&��Mu�"G ��;��G��`������g�8�t��&@7�U��-|���z�Ɠ��V�e��Ɉ�2�%+��?�������W�	K[$�X�ll�@
�mn(�.m���x��|/;���t�$�c�i�o��i��������Dhl�v=;;^����Ԋ���4��W���E�y�d�y6/qY'��;���:r��Q��C�e�Y�?Rtp��[QZ�r���KyX�X&�䟳������>?I~��af`>�W���)Ll����%�
���e�
d�0���xKgj�HxCu_�4lk�=bݺ���� Pފ��jȩ�L5���)����d�B���3�r�a�N�NQT���'O·ynx��(��Z�_���*Q�0�b�^�K"�.mMS��询a����o��(����aʭx7�,kf������w�D>,wRo�5� &[~��G_�q���ǎ�J#䋡O
X�r��_6Ӗg�15��(E��*Q�/Y�2� �ᾯ�r7I���"�	T�ya�x�%��s�4�:"m"k���.p��z��YB�:�{3�����嶾��vx��n#�J�J�k���:}-l�ɸ�J���VE��#9.v9�o�Vk���������[�d;������/��J�fhܼ���TlEW��`5Q��,����k�S/�aݑC�[�[�xRe�ݞ���IլA�o7,��G����k7����Z�����AM4֫�i./D��dQ�C�ə������~ט��r�L좽y�yQ6����C�"�o�i(fX��q�8w�"5T�Z�Pp��e{�RɅ��ᬞ/��������q��Ԇ�� ��|:�������5"�Xw��=�Q����M�'Y�@��
�G[H��g�d�A�wP�kZ]��g`q!�ϐ��^���\�3�f�怆�%/_��,�]���[X��<����8�����^����L�l��5!��AR�0������2湕6X�`a M��p(�ZA�j��ݿ����I��q�6F�Z 4�fw�4��;��D��)�=%ױ�U	��d�'�v�K�.hA��x
0�Ы���A&��V��!�Sa���x.`��c��8��N��)�R"��eƛ(��.f3= ��+!w��]�4,C�lL\�B��~�� �)W$L�0s �Z��//� ?W�J��u��f�$�ۊ˔U� �98�h�,� �g4�=� �g<��d�<Ў�O��
y� n���[��gk�oEڹL���u��: ��$|0.��w���/hT�M��9TF����ͅ�M�sWAQ����h�W�J-��/[�Ot������Ч�n$j$�'.e�$Tt��oW������a�U�����s�ߍ�ݡ��k�3�T��RG�? 773�Ua���c�p>���"�v��:�X�dg-w�Ɣ�ٙ9�x�
��\Ѽ@�@�c,�w\��:\c�4�7�cJf�P���v�Q��:,˵Ы<� �/�|���k''�N��j��kS0Q��D|�w32�.�i$Q��WZg�<[�9r�iΩ�Tat-�ROGI^�!x2i�0Ul|C�ۧ�u�x���S�^�L[j��NY��C��o�B8e��ǉ���{�̕�X [�F��c���zԵZ��H�mx�C�\iH�Y��o��j�p�����Y&�Nm���w5uޅ+�,>j9Dٝ�)ѻϡtn�'0K�"��EH�]]�K{Pv�2�{���q����!�j�mU�(�G�5�[E�bV����$�,7����ܩm�Q���Q���+��y`�[t/.0�U q-���}�`��br��H���uP��3��'�e�ۖ�q"�e����C��s���~:�3P��e
^ap�4��fQ��CG����%Za*Z��Ӑ�`�V�!D�%*��	ʿ�W�j��>��#��9�*6���)C,rz�,������x�r+�i���8�[ϒ�c�b�����Z�B8n�'z��j�tv�KO��ռ��v�Nz�g���R���j��.�.��>�@e��+�t��WR ���)䦞7��d��Ă��
�@Kr�(e�&al �mr;�М���!x�G#e"�#w�P���|<	4#�'�D$q����IMoI@J�Uy��ܷtx5� D�!��dĈ9xDfl�D���5��(T%�����1��+N_	cl}�<��x6��0<�oq���k�M"�'��m[?��"1�7�	3E�r�ׂ@���y��*�/��U¢�	����3��gt�����
���i;/�;�ğM'�W` ��ĀA(��X������s��0�_r�~Z�G��"N�=ﯾ��Պ~헻]�����t�!�(��A�7M�5�g�o�¦r�6^��J�_Yv�%c�[�8=�j��a�����궐�M{�*��f2�;��/ޟ`�1%�}En־:@�P%�B���-�^��33�F{���f$܇���5�
��%��t�6Q��K���/���E�{����qG���{�_FE8՜,��k#/\G��ǵ��j��尷c&��)(:���<���4S�P���<��	\��I;�Ţ��V��)jӂ}M�u�*��+�1J��&�| �=���M fՊJ�"N�j�X����#�L�6�4�ۖ͐9�������=�1��.���~�-����ӕ:PE��¡ <}�/ 
�'�+����U+�8y���1�?�����?��\�X�v4�iʤj��Xn���l�_�z؉O�(��(Wsjf63�<�A���x���+�*F���o��"��!��h��3��І�z]"]|��c}��i>U�"9��t.�j�5mx�	�����|�%G�-ử%�T��~ЭOӾ�Wi�w$��n(�����3~Fh�n�E�&��	��l0x�9䃚�����������K���M�A�u�k�N"�xb��F���=��냶��aD��v�,Zý�5��q�L�s����j��b�'��Z3N�/@�ѡ.2��99v���_�Ꞅ�2�{���;���S;l}�QXyv��ݳ��I�Ǫ� ?e����ǘ��^$5;��}���kI���$�f�|MP\�
g߬�cF>�g�=y\0'0����x�f��͉���Ԁ�y$���vd�B칦������|�^�Ɠ?�b��M?���A�UqS6�i9G�zk)pFb��*����\5@�����⏜S���ޘ�{��}A_j�,E�r���bm�>����'��G>�Ibf��l<���îW��̓�t`��6���#^ µx�;J�N��x$���(e�m���g���lo�nHc�ˠ����*�2�K��C�8�w���I�W��.�,V���v��|CI-����rL����=_9Q��j����7��\�QEΧm�ћ�>�O)�z1+,j���}8��:�4C�S���Rn��)nA[Qc)T���K��R.c���51�8�_�=EQ{SD_CF̜��SrB���yt�e���2C�_C���^�	�`\����Y�ᢖua���\��n�����������) C<NS��:y�Q�p�C�dZ^�7	~c�%ц>� �E�u_-�uOD��o���pVc1G�<���v�c<��@ߖ�գ#��cKir�A���#�`�|Q�/���;�ϥ�WAM�$��J�r}1��ؽR���ǖO6����II��a|�{:�Lo��˄`��A��:cN������6r�㐷G��P �'H�[.-�Whx=w���A�v�@_�G�|:^>�RP�TԊ�MYz��.���h��e11��3�{�����l�D����g`�筨e ��wfSL����pe�#>�gمs@������_RD����~ų̋�V`�a������F I �଒�1a���[ߛ�����Fc��Z5{���{$��"��l���]�^��vW�����*���	�n��z+���%HL���I�4�����কx�/Eix�P �^ɢl�mzc�%�-R��lӢ!n�q@���C��f��9�!sEzA���r��c(��w"&��L9���kݒ
�C��էHBq�O1��;\����	>�[/��A��'ֱ ��g�s\e~�ŀ�<����"���Ѿ�O����Ţ�g�j���t�5����(�r�Y�n��u�\�Y�+���#���ҽH~ȟ�\=�c�o�j�i���!����8O�)
6d0��Ά�T���
N�_5q�+������n���0(F�N0�,(�>`���C�2�*>s�k
�Wg��N��%LASr	5/��� ���$�_��B]�ZY�����!�I�i#84ӓ���b�Ȼ�.2&��0��U�s�V���c$��0���븋�QN��\����Zi��;�!?V_�z֕��_"$\&7O�n��@�����^��|��x�o�n� TJq��%����㞫مߣ�W}Щ�j܊�zA��%�a�
9z��Ok�E�F�T"Cdi�9Bw�ͬ�?�Z�v>&�d{	�Y@�SCo�*�٧K���s>����d��ǥC.v��"��q��8W&k�⢕��t��*�R�I��*kC����b��1�U��	����US=G��19#�'�B4a�a	r�K�^�g���]P�L�*kn<������DLbn7�@V�IzSe�Ҟ9�{\v��D����L�}1�qF�(*� �\�Fa�6X�b(3��@+"cWU��Zx�!�܁x9K�{&6��<<�����Q$�`�]S�b��,O}�!�*��-v�
�\2=�tW��>(^R�����Y���A�q�8���f����A����ph�' Iϕ��x5���̘��R����-���Z��ٓ��,�D�5f}q�6�5	�ټ�uM�Q���Cw��������F"�PLF��y�sB�}&+>m�VC�U7Dd�G>�dQrrP%��]��aY�K�E2�Q��N�db%�Uģ��7I��uJX�5+�L�9���[r:��s�׍&]�,��l�~�H�6�zߠ����%�D!t!sP�3ԣ&��N~��R��XB�g#~��h�Q{Z&0��6˛�_��}@��?�⡍ҟ��K&��9�e��R6��Y��?
.��
n�&���A�!K3��D���p��.�f>�*vr��1I�R�˅�α�L��L� �!6�%mJ!;|�y�gD�v�q�`��M�@~T��a�Ur
n��;�]eM��֜�r6�3S=#�iu��������ߨ*����D�Ƞ:6�j��Vy��2�%O��N��
=^��UA�"p�u@?��U����OeNIq�W*	J��+�{���{����;򿀜�)dW.�
CAܰǊu�ߨA㠘�FWAH��&�F���җ"Ub	Yc�*����%N*���*�D���,_.Z����L�r8�t�vG���=�LXI�RT����1fh�$�M�:��b�"����qP|��3kZHB�K9��چo�(��^��c��>ٔ�Wq|�a=LF�v/�]ì��	,�"�x�K�W,���N��a<��[�A_{��_
��A`��*�{0OoAXs�\��nG������hϩ�c�ŵY �.@��n�A�����w�it�e��������:o����r���㤂^}�"���x���\�+�ic��c��7����B*�#�CVr�&�X��"5�X3B��/㊠'���e�q�����̶ɺ�^�u���Tᤇ%��Bu�,��4f���Y�Ň��Q>��S������=`ѬI����~����P C$W˓!�t�򷌻(�9:��?re��,�9o��sިC����j�.$��̓����Wp�)g��;I�x�]/=��N�4zd�w>��<(QrX��&��q0�>U ���rz�_�/#l�#�m{�F*:Ja]�Ѻ�;���%��;
��Ҷ��0���.NEǣ�4�~t;���֧��ۆ�ۇ��ӢmC��@ �3q*��U�~?�y9XǱ��CF���"�K,J{|:���\�MZm+#�'Y���,u\yƄ�X
_�w^���]G��s�i���'ɞ�Ɩ�R���͑
�mg�l��n���hd��B�\6S&�F�~���tI���wm�]$�sj:�����pa ��U�hO��mpJbPB�Fh��يu�b)�Vf�C�M�Ms�T¡�i���eL 3*�G�!ϐ���J<�%2�<�
RJ��U��]�+>����_���I�ѭ&�pMֵJ����(T�i]��lo�(�a��F�h�����	�F���RX����t7�+����)��{:LⰢ�g/���){\<�l����	�[?����q�0����{e����pt�]��qc�I�S<"0At8�	1�
$W$�y�=K9be
�u�d'\���D���cyR���	�ǒ�+'�x�����V�A��O��m�a������9Kzq��S�Ɏ̭�t�4!�A�ofWH��H��a�'�/��\w�����u�f���BmK��N�9�� �&`]�{8U3_�Oy�ۡ3�r��}C���{p[	�f�SMu�:���q�m�!�����{˿�Y�Q�����i'��4yS	��R�$��H*��E�Xo\���~�'��%y* S��G�I&��-Ĥ��'}M:�#�g�ӑkWg V�B܇*x�+UK���~���Hlv��
�dAJ�zT�ՅjG��V���ԕ�R��l�FSo���hL����e��+��>�DQ�!�ېc��Oip��<x���w_ږm��|��=���Æ ��"�²XR�1aR�;�aV�ݶ(���K޳ѧw#���R	�Ŋ���/�2��7wdT6���!�A�8� T���G��TI����t��b;%�Y���Z�����ٙs��F>vuw�&x�	�5���ǿ�-�ӡ�7���֣,�	�B$����,�y$�Å��2�Ұ�w`��1ɠ�DR������A�{����<Vb}/��$�	U�bw譽��Ê����Z�)R u]`����
�ǳo���������$��iB�ze�ѕ��<eة�j���f���P�|��bJ�k�Eo	��k����e؍��G.��jNGQ�?5�س�^X�)��-T�0��Ϲ,_����4.Y���d���ZjܦI��y���V��������f%�v{EXP}<�K�[�T3�c4��"��Cf�� ����������l]����Ȅ�'�R?v�	>Ie�0^z����G��ٔtޜ�ܫ�!sE+��5��Q��L�p�H�V�٥��2T<\�5KO.{b/�;�皬k�E��J�33�X�<�2����O�J�A����Dm�U�+i �z7[AFgH���Չ�b�ӭ���>���3�*P2��"ĵ�����u�b��Uϋ%�V���q��FW`3h�_�Ը��@��X[P�o�W�tA��7���RC�#R���4Tʞ_~
�|�Z.�-m�l,��e�uJ��zu��[l�@_�)�[�N+2c��y�DPW��+{!�{��*8Q��yr�qJ��MĊ|b��`�X�7�e/^��Ty��T��:hf]��ڥ��9�����a���1z�;��B4{$+92���K����|nk���t�Ij� z�����H'��~8�њRN�@"Җ�H则EI¬@Z7l����?���|V:E��0�Z��۳���@�)��8{��9��f��*�O&�h����`xYP�ee���6��kT�8S�C�}�g~��W�_w���'�c�r����r~DE[
��ʎ1�p��w�K�rREb��Oc�\>��3�-H Yi'�����w�U���wE�Iس�%�&H���t�Ȧ��ˈ�n���e0�t��`WdC��`_3��\�J�M␠(]$0�Ҭ���J��<���5u�FR��	�����>�'�m[���V\:\~�|ܷ��@�<9�\�g���o�?�.����{�<�>��U+|EK��Ȃ�h+9��:�W��?f��0�ϰz믘2H.����n�Hz��(���I�y+i҇1��b��=�2G!��&���e, �K+�莹����0�1?�]��ȡ�ٕ�`�;�;���:n���X��	��b��T;'«}��,�=wC8zB���"���^��"�&Ёc�D��@e�H���AbӾ%K��L�D� ��.�t���#`�qJ�wu�$\�z/ׂZ,�2��TJ��%p�>~DT�,�gՔ�p��� �j�م��(qU��*�}s������3���x$��hPI7'�I�\������i�q�}j?�:V@*���AwӲ���ع��N�Q�;G��u�5)&��t/y�I��T�)�|���u�FT�ͦ"N�<�Mk�&��8�e��5pZ���z)#?�h���!&�~s�U�%�N3���s,&Ζ�g�C.n�/c>���˔]�L{ut��t��ڀZ%�CWL\W�ZbrYx�_r��Jފ��EV7<�&%gfp!\v/���b�o�h�X8+%`���5�S� �e&�&}�t���H����E���jnZ`m F,���"�J�W*D�ߙ��D���e,���Z}�S�"��H��C2�L0*k��М�����}b�G���c�u���ac@����Ǔ �jU�]�j�>W����B��|�� b/&�}m��`�[�a(�	�^�A��%r%A���e߁�������^]3}���}n'S����r�'�cW��J:�03�W�Ӱ�c�hm�M�ȇ�]�6veQ�i��y�h:�a����	gk�ҳ�������%�4�:1��:Ō�e���R29H��G$Ta�gj�)�@�{��s���60
�D��?7�Q�2.c��Ńf6� �ž����D5����	�C��XeGǈ�vQ��'i���_��oP`#���$�3z�R� I�ܿ�Gᢆt�0�S=F�ʃb��6A����aIEq�/��p@콢nP%$c�� Mz{��y��ĳ	��#�����G����I��CyY�]D5����_��|9Yq�?x}�h�ӊ��$�x�c��dڑ����4֌���J��q���;�Lo
�,t��<�FE�$�qi�t֢_p�2��woYܧN?���m��Vn툏���̰���Lܟ�$Y���m��d\�+�e�m��g+-//�C>+3S����
�˲��("�g�3� $��8>�7y}��O���g�J�� ^������U��B�0*�r�;��0�ސG2�Ot��7P�Y��gK���2�g��p��4@���ъBAh����c��Ai��z�B��R!�ޱB���/���wَUp=�?O&xe��2��:,N�{�,0J�����l�����>�(!������ϱ���������&�vó�������W-��ө�I@�2%�k���ʚ9��������՜��H�i�5=�j]9�2K�0I��A���=�Rux��-_�%}����_��v�IS|��Kc8t��mn��v�4��s��Gp}8����
w��Q��M�CYE���^�lISn|�Z���mg[�	Շf��Ϙ����QӅ������Y;Eƫ1uYK5qSL����S�D��Es�����������1�PwS+�����Qͺ%�'ܑ:vqɒ0��	:���z��;t3P0��]m�{�D1!;f�&Z��e�����>̑����6���
K���s��gZXwK5�!���L�����~n	�r%bw�4"�Oh͖ƒ_s�Z6��Ӱv�pŷ��X'�@����Ț�1j]1dh���}�_t��p?F��(�j�d�YOD�$��BKHB.<�F�K��Ȼ�|2M��궫�k�̌Fq����L��y_��K/H��)�8��P���M�#�ѓ#r�ީ��L
XٖNp�V�V�%�Rq?�o�OK�A���U�@ٕS�Po�*���>�ǻ&G���_�R�KZh��vc�S2b2Ց?tvO�5�G�ʵWR����oĔn8֊jW��z��3J��ݫ�*�@+���sw�zY��S%l庹��K$�VOA&o�y�ġ�R~�"$d(�lV��B���+/	�Ō���<>��Q�I�B6f��ȉ��Gu�\[�ŰV��!k�1���h#=颯�.���z5�C��>M�L���ꢁ�-��iޞe]F���	�R,kǥ� Z~�G�.H.q�
� x�59�$aaWw�
>��V4��o�1��(�K������S3���E/��E��6�r�m�F������Ŵj���P�2�T�^�^I�>y�Ƴ��ji��<s`�g�ҹ�X���=��h�`��ұ̦X������|�FQn�h��%��{�R�w��]�4n�t��oϟ$�N�mQַ*xl
B�o�?�e�=���"�S�OG�@#ߘ�ԗ�bTI����l�ϒ��³^��E�I�-oC����?����q}��/�#a��GE�؂���N��&��JU�r�-A�<Hmh&`�"�6��;|h�bMT���X�,Zl��{[9��]wXw����������.�d�p�D�el�����	�ǐ��Z#��;�Z(I�~B�q�*�)l[Vq|�w�3��ĉ�x��H8��?c�W�!3���D��W4\�<��	LXa�D
ҏCb� �9Qu]�4�CQz&i[�� N�a�T��%S2ܓ��LT��@�T^۟,��-��.R�����E/5U�d≃:?5Pu�Q�.�[����B8��g�n�c��)������ek�����+�k1�-4=F���]�������tD1) 7w� ��z%;��39Y�V �#aSˉ��t$���&:Ġ���c���̳k6Sی����P�Y�7i�O�~^Ga���z)+�̽��puU�"O8�kݎm?v�.w�2f��̈�u�S �^�$������X�u�S!��*���:�V9>-\���ioY����(��Rf [��.��>Ș�2}�኿.�F��z<Z��������"��b_��ma5��;�����:
��Z*���Xz	��N��NR�(���})ZyƤ��T����H�� x�tK�Wy�i�1�?\!+$l��6�C ��'1�h�c}v�RH�����q�(���Ϸ
��}�Hʁ�MT�VM���r+Y҅�>-2_W�<9	í����	Q�vY$�8�yT�
0W����a5�ͫ�D���S��X`�����-��M��?!��`i}���w�[dT�,��d(7����lރx�H�G� �E�&��M�*՝Ē��T�`�N{�+}�$	�+�Z�ݓ��9Ì���x>f��: s��;<'de��:ҹ������� ��o������K��"�Vz
vN��s���7K˧tc��jw�(ݗD��2�&�P�)���'�ho�)yq�QJ<�a��`�Pem�Pȓ�B&���I5$ �UƗD�,���>Q������-\V������3;]Ă+Ym�d�Y���H�5�'��E���s�-����42+A�����jr��Knj�Q�B�� �ZN����8돤~q��p�����	[�֠��{IY�/&Fd�}[h��(c�/I��N�e�8��J��l�բ�ٟ*��� !�R�+l�c����F��'0Xb��*���ھ#�5��ª��$I�@��O� NcM'G��]�JQe�������~�?�Wl�;�%`^aa��Z+�Y�v�}H��7h,*�1���`����G����a'm&�Z�[tȸn�[	����â�k>� 
8�ߦWdj��)��&6٩<3*��)\�7�fI�M>R���%�����~_A��}������!!F�=J?�4��	u4��M��g�ȏ7V��K���|A���\���2:R���Q����-��Q�!_���v��3Imqu�+E��?
�	hn �Ę����:&S��>�ν��6��������U��X%��v�khJ������>*�.��'Ӗt�������keJ��I3D��*�5�-�6'[ML�P��X�������vݡ������ݩ�n75d�(B���g�G�6�j|`]��u��&�m+�[�KzY䗜�4p��:�Ə;�_�d^��LNЦJn$I�Y���%�%���98�Ȥv�JxaO�M�Q�$�@�X�[�N����2ռv��mxA�����j@��:����׿�>q��Ea�a>�8T`��6w���Gg�e~ho}�J�0Q7�w����
WX��S�@G�]����#Z��|_^�.j�ڮ�@X�&O��FKI<�J�b1~�A�pm,�6&�F9zN�<|[�CO�a��@9����?��:�+$Z.23���JeΘ�����#������Ap>y�~���T,���4���ӿh��X�yˈ�j~f�k��9>�3����:�.[�����8�7�{D�D���p�r���$�Z24�:�����w����]������u!�1�Yw@��ɀ��@�kON�5��7|�k���bcab�����(c�xY�HM��m��!.�Sx�O��8	;��&��}n��9�{�� ����WT���`��#�W$���C+�����>��
��3y.��>�ˇ�JZ:�erx��]��� ۮ��E��ö��|͏6^��)Up(m�+��v�"#�7�[��r 1���RB*)�R��4��3�2�I����U�W��Z�r��M� bk�ez�E^R��dP�A�OE��!\���L�.Bz�] � 9������9�����l�0�2ɻ�}�S�eyG���\��T���^~�y��X��"=����v0�?�ym�M*�����k�&�� 'V�'��$�"MN��AC���vB*�|�t[���A���vg�8�xTt�}40W3�U��2�ZF�FLa�H qg�Av�)t)��2S��8�����V�j �k|��Z)��je�r��� 2��E�rE`����A'���0E�Q]vR��ɋ�2̷�&�W,���
�5�}����⊕��������#u9fK�F̻��p)Ӂ�=�/�яf^�Z��H�l�o��{�4u��������oְ�C���� ���{�|Du��AVm/�s_��/�˼���^K�@�_�K� �Rպ��s��쯙�[A�կl�+�"�y�0?Їt�J^-$�[�fUC�<9�Ґ�Rw��U���K?֧/Fѧ����W���}':�wR}|5 �$_�˩k=h�CӮ�q:��OlIxSO�]���R]�Ƽ8����F��A
����)N���]�U��tԘ }s��wr�@� ���Q_1��W�S���������F��Ċ�zٚ_��m_���ZT�G�ם$ώ0U���]u=����mda,�}_����$.���V�a�K.iɈj��ǐ�@U�v ^�H��,�7�
N]�eߑcwK���L>3=����j�{�qT��bM�rr>�B�;������VWM��2��^cF�v�MD�C�ʡwR�EI5CV*�!%�C���(_-�]�,ܪ`��q�W�[&$�&�L��34��B���(��� )��rlZV����|9M'���Z1��ӵ��r�תZ��~~]�d�O|�eS�M6C���,g��
��E5Ys�
<�w͖�u+�eA�+�Ӣ�K_'�ś�����qF$4��|�X���ӗ�ߩ�?V?I��ָ����U�&
�|�k*�>We&�9A;HE��y�t��D��;��Y>�����~�l�u������3�^��{���r�Z_R�^UtY��u=�w>�i�T�$�������:C��ր��ě�3l�a�$s�4�($7Í�q����e�{���k����41��h�����lyj�U��$�J#�|�a�+�w0�"�״f���*_i�����K�!${<p}I�� <����bu���mf������z�Q�.��O���=�$��4����uݵἠ�����x̫ ��y��/q�I�QYJ���~ �}u���V
�Dtf���pz̝c��_��[�:`������l��"�xF{�J$�}͟.�e"��N�v3�9���
�R��=c��	w��2�vR�7��_�>�r]�+F�>���(�Ť��j�Ps���2R]�r���U�V��1��A?
�G��^E'�)���Z�Ynaww�]Qk���P��>���A�y��pn$���� Q�>JL�p�-s��,W��ƴqc�}��	���eu�.���FhήX�7�_�*V1 ,$��	�v ���ז	�`N]0
��6we(۴!4�z��iI�}��t6�)�M�*t<}2�1�K�h�(x�s�,���w��P�%WY���@E�xߓ�}:� �>kg%���ܑ��6�k����������S(����#HO���A5(a�LSl���(���R�������&���}����C�7�2�X۷�����>Eu����rr�BGH+�o[����G�àW�
c��lzS�d��;b��N��?�b�H��A���G%�ubz_!E&��06��d%�Y�m��`�̒��/��eWbu5�@��JW��V ���:��Q��ٟ4t�Aѕ�d��AiJ���	kpTۄ�U����ږڷ@��d_s�j��l�z��#��I��8:r"ُteF.�9%�@�\��� 6�/��(�פy.��_��ѳfٕy��B��P]=�Z�n��}pq�Qʺ�m9�^bC��f��g)��0��}��ʜ����+nӊϴ�6�tΙW���oF��!���X�~�'�S�ܽ�F���A��U��h��<���HUE/CDu@ȁ��y9:�:��EѢE�^��8a�'��	Ƈ%�0��%N����h9��\�]���1�>G�'1�V˽�X�n&����`�:6�xRP���(�n��3DAݯ�O"�۰�ui=	���r�()���`)��'k>��?%�Fc�"N˱�6�Ȏ�bo?�����8����ɾ�V�)�L�>�cHY/п��0<*��z\W�?�;��X�u��Q��;�+��7��&_M�L�b5���;v��C�r&/��X�C�q��ޗS�,>�Q0���rb�װ����{s�J&e~�P�0�gИ'�Re�P� m� U����B!��a�@��(�#���Od4�3�@gU�/�F�{u�$���`
%��>
Ϩ)�#���8��\e}�F��v�3�]E|i�v�gr��Q���&�iX�1�W��#-�5�#�D�0{o~�ie�y��N�4ґN������b��+��!��2�/1�476zfR�V�惈*P��ȿ}�Ĳ��풞�ء��-"7\��O��t�H���kS����˔ÍU�\Y
*��+���Qڙ�<G4�L!�~U8i 3�X���� LsCh���[D���%�����u�bs����F�
�~_�]`Y��n+��R|�vk��7B�
vAI4��?y~r�Ș�l�p����Nϩ��#�F
aT�q��e��z��Ģ8��(F�;Q�K��z�'�)韻%%Pa�\�"��E�I�\�4g��my��=����<`�j^e����;��d]����O�hpJ�,����0�0"K����u!����ӽ?�vg�Fi�(�:Qz������/h����-]Kh~1��ӮJ���~M��u) ׎{��Z^E&ؠ(Dmc�o%�!{����漱�=�MU��b��6̀e�<��X�P?H{3���/�F�G.ф�/�4�^�:Y�k�?���=��/���Tw����B��;-8\U�F������:I�l�"��>��S�|��P!�
����x�N�^\� �v�q�B�L���@,�O���;[���0��Dq�&[=0ml�Uڅu�b1 f-N�B�O��l��D�����֊q��.s�o�g�%8��v��k�7ݡ;�G����KA�"\�].`�U�^�b��%�:��3�<�u7���ڠT"H�to����ı&)Z�{y\=&�9�(��ꀫ����Q�Gs�#�k_�8w>�5�7�� �)�10�d ��z#�<��S7�e��z+�oSeC 9xE�z�%�rQs9�xu+��#����M;m(�%+�f�U@>��c��Μ�CyG��C�wݒ��eQB;C���A@H��=���Ii�o)��!Hyy�q���5\��LF��R�Hux�DL[���qrV��D��w�j�2�_�B$<����njQ����qiEwZ�T�H�!^VD�J"յ�b�7��'KG����:B�|tn�?�
�m|\�؏��f@M'W(�f�K�4*��aZ�Z�eÿ��Qi5���(ΎLF{_��YX�.�p�+����5Ip��}�!.4�Z����N�<���|�����Yg� 	X2c(�_`��C�H����O�\FsB!�H��|(vf�{��hjƺf�����Q�Ω���ֲMm[i�i� ?5*�|j3s��������p_h�ê����:�gQ���$y���F��>��mxŠ�ŕ�"ɜ�n��~�z,���{�L��$���m<��IM<]����Ls�d=L�I�:ihA�33E���}�.��xAC~*�����צ@T�C��ӔX`���O���_��洤ww��)ݨ��Af,d-V�¶��񄕖qP,e��d�L��hl@d�4�E:)������㖣a��/��>�O����E��^r�;B��Y�	���u�o2�+3b.��-��_WM�tg1��V��A���vh�Oc��Y6�������f�<�����0s���'\��DR������6]�`���(�1.�Aф�#piZ�
}��*t�d�OxU�,�WHV�t�䓪��wwo;b��[Œ������L@M�����a�S{q��Ur��Ib]h�p�M5��Vr�U�{���S�JX~�|p��#K<��ߦ�c	&.O��*V�u�� �zH��<t�Q�C7jA�����W�a~B��5a��/})�2��~�U0։�{�,�*�����}��gb+S�:	�b��u�Si��P��xdM�aK�+ԥ�b�hd�Bg`#z�K(�9
h"����g��.�7+*�)�ϑ�|tz�)�2쾡�F�av�yi��P��.k�����D��f��p^1���.�,	.-��I�ئb
�?����wd�Ҏ�'k�CeƲ�C�jgW��ÞW^��}w���9�# gh���s�6�����z��I��*�dƤ�K�3/�����Y���;t� ���\�o|-o��f�)��0��ѹv���H�xڤ�;˪߂�J���]��L�2�VO�'Ӧo�<G���`D.Ĺ�����
ЦS��",�nR'�^B�v�?!D A�)���ΚSr攐�J�&��gG3��e���LE��B���s�Й٫�>�ljͺ$&-���I#�t���6p~��pܫ�`��:vI�u;ć7�.�
��e*7��j*�J/���{+����u43~,On�@�=M��'��S��+��?)O�w����;D�u0sA�Aۿmb����D�hPo��iѰ}�mwt�P��+�v���+�^m��Z��)]�w�\�"�: f��p���-�'��1��7x�r�S�Z��xv��.��oO�RQ�s����������j�� ���S4�[8�8�2����6_$����p!��V*���B^���IW�H$��ݡp���_6��c5�D��p�b�8-���i���v�zԜ�ۣ��0�E-����\=X�����ĩ��4����� �ݍ�\p��ו����/�)D���p�3a���LE_�L/�@��^9�Wp后��v�<�k?Q�h0
����/��4���a�������dJr���D26����,�&�$�ե�'w��{����B���?|<.aS�" ��}��.�{Iy�M��������}�%�`�#t��7
/�ĳ�W\Ԩ&���9C�TΝ_#F��h\}�Lo�Z��^�(���c�����K�`e����?�P���¡�Ln#�?5�׍ $�f�5�'5{>p�rQ
'�oSn.���8a����O��*��>�a��`E�Z&Vb����~��n�h.<�o90�ߖ�-��,gY.���ᗄQC#$��2���L����+t�&���S۰��"4�}�Bցb�U��q��T�@��C�aN���$��ܺm��x�M�\�&�C.�jgW&uR�_���*�`�s~^����7�$�|���K�������G��o����"�$��>C�����`R�.%�c8a�5no6+�b��k���-�~����4�Z���o�WД�L��Q���p�#	��&�����Rx}�K6^��#��!��-���7߻9��-�+D�hY�<�=sn�咈��C� Im�/���u��t�;�F����Ҋ��9�q�O����\;sd����6��#ǽ ���z!~��GT^1�7�&���9}��Or����  ���P�V��ȓ����� �!M(ΈI�K%m�T�Q�]�)���#�����l��:�=����,
�^G���2cqJ�@���;���{�&�&A�F��j��Ї^�ݯ���jmu)/V=��3nf�6=r>���,F�%�o���H��J�"�����g}ب��N��D�qt��`��eKcV�d؅�bM�-����>+]6��x��_�7���y�}B��1d�/��ɺ�u?�J����S��Ѓ�V�6׼��$��~�k��GL�SL��b,D�^��D�{�p��9�N�ʋ�G%\Z��~I�x�3�ږH�H���ġ_rM�y���w�)vd�1O�ؑ`�ElMg�1�Ĭ܉��g�;�i`n9s�9�����E���Jp�{�$����Z�zOe@�~[�*�����BML6�MfU�up� �횄r���-V�HrV�jǼ�c^��%2����lm�Z�r�{x-&��⦱p�$�b	��f����]yC판�6��������;e���u&NS!�;�>{^#i^LE��Y��G��E�_K֘L!��,+�/�9rH����s���1�����'f�H��y�U�E����cԘ$�ɶgRV���G�l��H�������c��D~�C�>���Q���p�)�y���~��l1EA��:tܗX,N�ޱ�kh�~��Βu^�C��|p���u��炼��a]6v�њ�N�C�U�]h���NCTZS�T�`�rj���c/�،�)��2�O�q��G��X�_���]:��a�=�J�1C!䊽N�7���직�8��( �EX�В`�a^qrPJ��w�MGHX�^^`�-8Ir�Bh'�8�~Wy��dab��6֩��=�@zg��E���j��<E�u�i~ks81q�� &I<'4���L\LC;L]y�>=����Iy�͝@Ts��֠L�)�e�2b:�M4p|˜0�"�J^&:So��&�^��丿̉�����{�9t�WsJ/�[�f�Du��ٸ�$���F�N�Mm�ﱾ]������xx6/f��a���X�π��rJF��-���B�ޮ`�rc{<��������/��֪����s,:���K��u,>� �?[c�|�6��A��`פʐ�ȸ���
]I~\��G��֌�UGK�[ � �i���J�w�yV��8԰`�8a��t(n�k�L���j蒕�j�|]l�om90��O�˦���.�6]}�u�J�a*VnW�a��������8-y]$RaK�1j����ӌ���=�.Kð�\���#�Ѻ���1�����O���A�Nǎ?]^Ӣ�o��]wo1ՉS����N�<½�� �2�͵�.]����o^��Y��m08�Y�fǡ�x�gq��"�V2{#u<���<<+pfe���ph\f��ɦ�$�%��}R�h�3;2��������:�q}���+�%ڵSv��m8�tU�� �߮���/l���I|����q�	�v4�#^}��=�3Y�F�Qm"�qT~��	jJ?-/����(��⊫@�[��������q`#p��W�n-��J��%�N�<+(Qز=��񠓕F/'���P�j�I��ż��v�i��i��N(5o�<\!��ԲL��09�ݥ�3��-�agV���zaM�װ���j���T�_����87%x�����s	����c��M�Fj���3E�O���ɏ=s���kv>���B[���#tW&ᐰ~�RΞ^��F�j�0�> Y*6'��=�L�@4�W���q��F��@uw����� �m\&�)��~��K��#B1?�]��le3"�B�HU!tP(/��tD�����?K��w7>b��P�\��]��Lm�����.�!j���,
��� �n: ��#8Ɍv;�"��C�Ϝ����ہlR��B���y���vЉ�����3�sOL?B�_p����2]�]��6�$K�(�Qy���r�$�d/����� �#�&�y�K�o5ktP�OD�1d���+˽SQ?�pa����qw#|h����U�g�u=ƨM��1�L5wm��,j���vj�C~Ys9q�e�cu0������]2���_:���}e���Urp�2�� '��z�������9�9!��M�Gn�A�]i��sA:��r�<fC����5p�įvǸ��{��[�ҌmR��6�~��YgW'V�W_��k$1�!���[+�?�������9퓵���1&�pD�G�shN��ER�T�Nn�G��1ɋB���>�-AŌQ�Jچ䶞��m1)�}�4A��
���q��k�c6� Ts�I��.���M?��u�k���d
��֧z��
޸�n�zv]zqx�~��K��M[�����һS��tff7K�J���js���\Oˡ=fvi�	� ������R+Q��T�M�uzM���%/��W��.���U�x�1J��TK�ޭ<cƎ��p���N�m@���b���5����n�+rV<N�����!k	$�������9> �\�s;<һ�RHe�JG��b�������q��D�O���\�gg�������NZ�σ�w����[׿۠�CE.����O. sqz�WL�9������&����1�FxS%Ѱ�-"�x�|#a�Ώ$�ˋ.�X���� 7�)���
w��Ʒ��z�^�7��3�>����Am�_>u����0���N�Q}$����óD�Q� O4���J�e�?F�Jv��N�{�M!J�l��5�8P��
��It�[+"|}�k.��_h��<=5%2�L�.a��r<�9?p�a�0��0"*5=�=�L�1��;c;H*l����R&n�$�B�{Q��\<�����><W��Uy<�d*�}M�|���5�ौ��ƢnӒJ~Z�.�,�Qd��CKbX������:��:d�C lM]�wv�ܾ���!OHr�0���ODj����<��q0}�p���G~[��e�����`�D{Y�ĺLHFE�=���No��V���p�	�or�M�z�D'!�hS���m���8�vѦO�[�pZ#�H�JJiLx�^M�|��E�$Zos'u'����H���c����~<7yöVݴ���N^��«�lf*$�a�@͖�&_����,UX��b� @�i�HܖI��Ǝ�"+H�c��\_EWoy�)�`KE_|!b_�+Wn�s���b�`m���'�+r�r�p-���Ţi	��R
���`D$w���w�l�Qyfn�۹jF��"�?h�����?��4ƸOz��4uvŎ�3�6FI���I��x��9	�o�RU����(^�"��B�i�;\��+ ��p�o���(�20T%�T�u�6U�S�b�>zLř��	N��2�q�\q2D�~����c�*����z%��Oo�:#Sn��ݔp���p���8��6.�=�{lשm�g���.\{K���s��;� �8{�W�|-H$C?��G!�HC0ic��Q�(Ѩ���o�PU״`���PT��[v�Xu�B~�h/;o�#���@����'ܲ���j�v�ob=�c��0G���XɣP~��������.��<�-�q�ܾHlxt*��S-F�m��
�W��c)b��҉��~��ţ�ͬ_�NFp~�V/qcf�Å����b�钋k�65��	*1�0�`���l�T�f���H�8�Ȁ��{yĵ����mr^8����ɲCa{؆P�{�&�}�֊��x��=�FEgԝR���$�e����`�)�H����_�-�s(;�X?���+�1_R)�YUP�1' ���.�`w���}�*N�$H+�_����p0H�]��]��.cܵԀ���!E(ɷE;�,Md�����XL�>jI�ӷ�C"�*���m?4�tCG�fg-�k��rE+.��1M�f�9��c����C�6C�{�q������)��>�32�JoDrjT��!?��߷ZbC��
�G��)��Dh��_�k"n��ݴ��N���
m�=�F�x}�A�_<�`&]x�{�m)�mΥ�ᵄ8]k^�8� ��lp�x��Ǘ�
�宆�X$�f����Q��g�#bvdR�/�������[���C��|��z�?-0�hȌ�A���4{��B�.t�N4Y����9��+�
����WAP�
6�@��	�[	<�
l��C��-���[�#�ؕ㊓]�{w��|�@z%Y��@��ĖW��2Y1�,�9��򖜘��e��,��F��'��ST�w�f0g�w�ٵ�Bㄔ`��n�&G���,�����*pƞ��qݣ��5���w%{f��Ɖ1�W\���&|s5&EYx�fW�*հ{,�
��"�h��]��Ѥ�N���	W)��H{�F��x���zD�%��8�E^FG-ǔ��	F���j���dq.�#�d{��Ƒ�!->����c��V_�mOa���;"y9�Zy��L*����Z0e_8A�P.��as����S�m�|�0d��������wpm���H�:�V��<�<�yW����'��%���C)�q�[��NS��q�<��f����L\����?V����q8K��P�
�[X��(?�`�����+�VͬgN�]۝�Q�j;��%�G(쾰��*l�I ����]0�<�ƄL�+�ՙ@v�&*{���P!���z��OF�|�o {�k��d�>�l��]3�eڸN��=b�K��&�1�����A���k�A�z~�����Wș�Ʌ�=�ð�q�2N��>F������ف Qf���F���O�����L�b�0��4 hc���cU����d�� �`��9�i��yÁ0P���7~�'2�挡c�?v�9�$�gO�A�S��w5��4�2��(Z^3m�s��3�Z/�:_��uE�٦ ����+D�)]�>Wƴ�ud�af��� H�5U��*��I�cҷ1<��������� :/�M����d��X9ZJ�q�dR1#�2&8̉r�T�q=�{SM����m��ݗ{��VDm�������?���(�]�W���F�'�5VH�7��(�OkR�L(�c⪶׼�
���27&�1�b��#I/��O��;�ޒ�7����fb}��vQ�~�^� ���<�0�W9���>[��b(v8����7���:��q��V{��L�E?��cn�	���xs��Y�����@�N,��5?OE�
S���,���e3���^7�}+�l������&�Y�Ւ��hV	�8t��[��p�c��<��|�kK�������vTyb�w�a�(�;x1��� |Mg��TƐ��X3ݫ�����V�U���\7�JWR�n;T���:H8W�2/�=��1�8g<�t"�&7����z��d��C oCSj�n;�Փ��ʇf�By�����������հ!!��%>�K�F�ǈR����YW�@bt^d�N0P��͇ڈ�G���=z����O�_0D�A*����z@��h\k嗪xa�WR�40�(�t�Su�+�b
�;�fi��W�(���s�F����b16B�L=��m"}#C���9�/�o��,�E1�ɺV7�Yoc�5�7�,��9,�wE�� ?'�3��y<�_����ɫ8WR���̯��Ԏ똹���RӔ_U��zc��W�8�ϲBO:��ɂU�"vu��o�0�k�0;����@g�3׃�	�-e��P\�V���PVJg^���B�B����`�v\r-tբ��L7�1��`U9�y�K�V=8�aV�02�����;�W��j����%�|�֜eV���${�~ yz��L1��!�w��N��@>���M����9��.�DM������"�p�2��|\�?��J��%g����٣���R��~��OJ�oKy0\��PR��@����1������"&"��d��1��3r��b�����I&�yeK�)} X����E��?m"Nb��a�B�������KF:aj�)��7�Nb������%�ː�ꍕ���D�i¼M�E��֖"Nh4�TO�-�_���;� ^*W��FѨ��PJHA���K��dN`����r�|��n���X|D�w$�H|�o�/.�i���9g�g�B���^�i� +�@����Z��Ҁj.�J�C���I5P��d8��x�����*Wl$�g�4y��j$�����7M�6((o���*��x�j���j1cvr�G�R����vl\�44������}�~�2"�ʽu,�KuF��+��4zl,�n�#�P��8�����fҖ�����E��C��� Ӱg؀א���k	�@kA:Tvb��p���&J1�+�cGi'$*���q��S&1�Xm��A�����x����|ysF�8 dj�A�(�g'&>�Tt�B&)��k	�q�K`�k��ǲǷ�jZ��$�Gi.�&
h�:�����P�-���h=&��-,�{@s4Cx��:P�7��)�2B
�
v%���Η�WM��e�
fg"��gVsKg��ՠ	t*��[��!�����m��� �F���V����j�ҁ ӏ�5~+�#Ҭڷ�gADP����$��Ǯ��[��Nۥ�J�)��2�en� Jde#�}s��nx�Kϥ�t���:�-m��� ����ht:@��\ͫ�'�6�"�#n�rSƆ�Wɒ�5� ?��\�'ɋ��߅6aŝu�s0f�������b�Put���Ϯ������0��ȭ@G
|HX�8�|�f����G�N G=eF���2ݣ_��9&%v�Gi�`�#(z�d�H��C�	;�_@�`"��5?�L\��s��t��N�ς�:�x����B���E�p�t�6'�?j5��t���k�$􂅆{`t��D����4]LA�,�p�,4�%\i�b��ʤB���Z�r���o%|��W��B���M��Y��͠\��y!�	�
{_ �������Mx�+(�(ň�%F,��(
�"Q���P��s&�Hs{����V��6YH����U���su�f6��������|�sH2NO�8��D���	�x���>1��3��zJ(67��S�L��.���e�"hgڱ��ݑș�-TS�3&�% �e���Q7���ѸHo���ݮ��"��cr��ϣ@3�T5ZZ��D��CtM翯�j�p�k�������Ĵ|cR�?����
��'[5d7�s/Nw��L8~E��NI=h~a��9�"O��(�j�F
f�^[Է�o�0y���R�x�[Z�c�\�T��x7�,i�����#�T;z��4�6"@��4>�Aj�B3ƜƂ9�d�ڊB��.�c���NH����m���}X�q/�Vɽ��3�v��W3��?5�ڑ��Ks��t\�4Q���A����R�+>�8f�le�}0֩�_� ���,�O� ��g�o0S�۳Ƣ,3����{҅�Z�@��BC�ø}T'U=&b�� �n�Fy2[��x��>wa$�OAg�_�:�w���i��s�iy�KR���b훿s����K�C�i.��%�ͩ'W�����׏M��T�;���-HG�E�"�v��O:(f����U���yB�{^���N���U���ZN���~���:qO����q���`'ىo(k��4M_�l���oP�ϗ4��_�̌�&��٦�F�ƚ����5��^��^@w�i������.u�ߨ-K(Xl>���C�"����J��J��fV���c���{{���/H�O"!��K��j��ʗ��dߥ.)Вk6�~���0;�V�qǟ:;�ࡡ_{�vkU�I�
x������Ɂ�/���hk��9��X�'u*e%�.ͳ��Û��5��T3��F�kֲ�e�9V��;8�XBTa���FQWE%������p>���a��շ@p7g��:-���'�F�-߬87�#�T ]���&4�SҾK���l�Np������M���./��`ᇘ�n�����X�ܲ���X>������<�!�x0X��I �)��2:ޫ�Wm�5��Z���F�%Fk(X�x(��~)�vG!�6V���ӽ7�t�[I��?�` ъT"Q���5c{s�?�lj�ٛ���[*%��#\�]�}f��� (�ua�,	����Eî�`B6$��f?�լ��]��P~M�Ԓ�,O�I�W&;}���5
��ԝJz/#:w_�G��$�h�E+���wa��T>��<Eި����`�&U�W���^% ��O,�	LAS�#����]������A,Z�U�ŰO�I�?�6łÏí�����\<�xU	�ų��^�}eD�99N��U"#4�`A.��!�����M�aL%'���#�d���M�F���WO�&oh� H ���]�
��X��{��1�O�/0�"r|�Yԙ&�м:K�()|�Ӽm$�N��Q�Y={�is�]1Qc�'�{�{���I<�z�=���y�o.���St�W̶��7�eU���e2��[5��R?\�3&�� �;����GbV�8�':�#w���`���A}� ,��9��^������Nu ��F2��q��s�f�z��Qr�7�	��ٯ&n�JhM��<�qK��t篥\ly��#�ڋ͖�9��D[�WH0��)D��=�[�t�]������Y���wZ�����G}�3��YQ�I��#���cws`5�ND�9�'UH��>�jW��Y�^QPB�W@��J�Ak6���u��P���D��/��X'����<'�$�	�f�u���B>X��X��Ș9��5W��r���zs�-�&�g���J����0ȇ<3#�b�������7mI��U����e��ϒDE�q &Gt��hǽf��mȹ���搌�~kg��}�����8�'C�O�G(y��j4u�G4p�g�I�+X]�6�I��U��?/.~D> Ԓ�!tO�F��~X���x���́��}]����"#��y�
�kFqi�����q�_���S�L���|����V�Mt@�AX��SL�X����C�iN
c����l:Ʊ�~��7xM��	Mx,n������kɣ�ahF�kPbXN�./^�t�O�)~U��}t�Ft�tr�!�7:��R�0=��G��NKh�+	&m4�@����ˈ��a��f��:4t��:+� r���m�|P���#S�%�
�1}�{��W���-�D����*H7��`����Q%�J�A�jy� Y�QZlw	�܅�����x�n�Q�se�B�Q��� �J�7�x�07b��.�dy�zњl@�[M�q�����oo��ʺ��O�8d���ǅ+3Ma����uK݀7Q�d2�����=��M�ݼSi�O &�}���ߗo� oa�{�߇�c��y�o�o�"ĩA������6ci��]�<��\�U�o����8J������~����ވ{����gi������֎CG����cR�6
E��~�Lg/�'pV�+x�o/ ��y��Z%9���~�g��M\L������s�K�B�Na��3;u���{��+�-
�s�)�VQ8$��״�l��s�c�׿Z��O�]�Ģ��*+�W��Η��]���˻��4��g#��j�6���j�s0K/\@�p�S ����)��5 �����(�0�A}����x�d^)�ϳ汊�B�IZi(Hd��E�O�2�O�X��%���D�Iv/�O��B�tw2����#8w��ި�dţ�M������Iay�0�%��1%��ؑ���v:D�!������C�%�m�u�<e<,��cm�$|f��6�]<��c��چMw�b�UK���ǿ2$�f�687=��F�
�R�V�����^WX�ĘC�Q%Ѥ��܅=���D�G|��A6���}��_��G�/#<Ρ\�A�&�#!V�=����E�"�s��eI�3m��^ާ���q�	��
�T>&[8�a��v4��sm�UH��]����+�3��q#��}Pd
�N���T��k�� ��.�{���\9�X��Ʉ�XQ���~�=ց�{$����%_��uo�8Z4���@�䎦��О��. VT��kV�ģ�rw9��� #IH�oy�f,��9���l`R|�Ϳa�{�-��F�q�F3��<�'Z-Q �\����}e����X
�����R��
G�WGϫf�~Ct��ڥw�Yh��!{�&xK���E�9�xr�C武�a�\�U~'�|ˑ�t�F�5'�(7�ZÜ[69Q����Qfy���x_�NEU���|/�E�E���j\�XDh�+d�DkO�}������X�ء�X?J�J�#Y#������G�1&C4uzH�O���}���3�V���d���gmt�wV�|'�!��&I�<2��Q�3o{�Q�Q�ۼ�)�c��6���8��ԉ�|�TaE$���K�<.����VS�Oѳ�z�����IԌ��RV��/�����}X�ۿ�5ZUE�+}�6�LNt�!i�>���k���@d��?"�M�!��b7�kV�.fJ~Lǫ΀̈-��5Te�;�f8���[7��Z#��FFs��0#�Y�%1�P�C��h��GlFr!CUT"�i�i���穲>�}i����%S�o�3���� �>!x�Hǂ�9����ܨ��럸 �y�I>��sL���O@�N�Wo�|2*dz�E>�{'� ���J�}g�`P#���w+���^ee �`���n/�6���C!!�r���!6-����̡��+
/�	%����y��Ya��}v|��\HU:,E��kx�E��)� a��&��Pzߛ~E�6{��}/�0�s;��W7��H�z��Ε�=.�w�q{E��R̗� ��	�?;,`�9Po�:�h�d��H)��뜒M�S5GY�D�!�����MMN|�d���e;�Pw���i�[Qi�21���2[�]O��Rk����G�W;Wm8�O4�HQ[�\؄�a:A�.��
5�'�(��v�.�j���#�� (�_�mb���w�����E�R�w*�7�[���[�Z�ҋ>�.��{~�d�R ��u�׮e���.��f]�B����ҏ��R�3���)�L8i0IP�\�m�(H��`�mi��'�+���<y�w!�S�{l�nc%e)]�w��*t��ȴ)�n5K"ާ���PAIV�5�eUv��r(���&d(�q'v�y���� �H܊x�T4�?�!]���G����ю⍩�UͿ��9�����.���$�����kȿ���?�@kb�r�Xpr�4�}Aĝ����åt⿾hj�ۇ�'*����co��-]����� �0��]<έ��.eE|#���@��;��Yp�M����M�l���Ƃ�!��6z:�B-�e����gEv}GI�~?�X�	��{����$VڶջF��xҡ���}�냵�u��棺�8�ݷ%j�|�����#�u;�XHT��_f3@u���nG4���D*�&�rW�(�S���huupi@-�\Ҙc4J�)J�\�e0,z������j�Q���[�43،�>�avaa�Q�b"qַ��r����㦧ܸ�)�Y�ݺ�s@���\NZS�@�]�����Y�0إ�ˀM��ج	EH����:X�7�������@�}{��
�њ(}��>�=&�g�-�Q�7�@<�_���A���m9��@��ie�
�g��c��T�yi���4�ch��`n����H��*-�%�@��t&��btS� ЌБ98��Q��d�����{Y+s#m*b�x�q���)�\��z+����F-��nn.	(�S�dH�)[��t;HM�	���j?���=���Q0%M6�d� &�E�}uϟ���������S)��`�ޭ�j�*��+t�A1��,�a+��qW���Ǫ�>.������>]��\�6�į��$�O�"��C ��ĒuP���tK��K�����B�ސ�HK����]Eqx���8�胷T �-�e��ٛP�-�x~�{�J���B��,N�Izj>��>����Z�j��������{�uUq�G��JKIAY�wN��D�}_��eS7�vS<7�ƊD���|��n~2$ὓ�G�b1?,(G4�������p�|%��S7&���źnRKE���ő���Ue�|���{����(�Z�i�t��L1���(�d�h7.�l����4Z��9��y�8���-Ǳ|��ufW�$�s
�<�xЏc��#n�in�L���� �ڵ�?�LV����8�F�Ձ�����E�ݼ��uV�v�_~d�{�e����B�h��>�O�
q���~��CU($���0���	ρ�:ʌe)@H�`�
N�#̡q����NL3v!���pn��6��raJy������)ŕ��{��k��p�Te��X��c���r+������>?Z��yi2����dѽS�.JS<?Qqq+�|X=�G�a�k��r)ު��!|Br����.Lz_5f�~ږ���Q����Z}P�!�c��b^��RgsYM��K��O���j�z:��$a-��$��F��D�S�6��I�M֬b���Э�"�U��ZS�A���w)J��ֿ8Q�J�֪���}�d�6���J`��pC%��H�+�B@�AS���b�2��Gm��
l���;G�C�+�o|J�*-�K�ќ:I��p3��8�#��D6sD�Ѷ)��e����Ú�Dm��J�-��α+*]K���rt��(,I�?����I<�y��*�����³��p��@N��E����6~�I�]nD�y^�?�V��ʻMdO�=x��Z��Y�����nwX�8��&�3���
�'Y�t ��ӎ=�rCxc�sQ�q'�*Ĉ��S�>�
��=F����/�4�D��bw$�\��Zz4��L%����d��P"����>�U� ]��4�#�7VFh��f����I�ƪ�>Le�]4��*?�\鉎=_*�ýQ'z�a�G����%#�<���;8/�qX���X(N���h�v�+D>�_�6��!X^�n����x�|0S7��u1$l54;-��K�V:83�� Nی�,��u�6�9������x�7����Yk5f��v�+>�o��*S�m(�O�5~��1>�g�r��[�oPJ�@!}.�s�+L��!.��)'�����y=�0柛 �m�����[$5�L������yU�fAB(�rl�Q�|�3!l�2;$�bkaRp�v9��ii��O
�5��cJ�W-���k�e�iP�\˩�ǖ3<;YP/~͘�q���s����r\.�]��+�-KL<�n�ɧw>�&����vO�i��d�g8�s��=��p{n�j�%0��a�Y �!��B֓#���s��S	�|�����ML�2���ݟ>~��0J$Ռ���-ט�y��i��Hp��AOM���R.h��;��G@�]�v��)�\*���yfw��.��XB �����g��Q�	��w��:��횺�^^)�o��⼌�{O1]O\��?���_B��Ť�~�R	�s�ǿAD���A&���S)���5/5�|P����8t�Lz�s.�r%���6�9"��b֧u���2�|޿��yQU���k=zL}�;��8cϟ���
��S��_@����}�#Q��D��+����]Ss���E�|55��;2c�~*�.�5�5�]������9�P��7��g�'�Jd�P�����p���N�WKV7�xZ$T���'??5? �8b�k�b�[I(f	P2�F��g~m�3k�/Dn\{�J�����<�Ki�iA8^�uym��q2���������We����Х'M���q�V�F��	ck�)l �� �-�_���<#sǀv�yXX �� /���]=Y�j:غ�U�I�+4GW�&7�KcI�R��ݶ/U q��#h����]�൑�MI�"��U)V-���;%���.2�%wz��-Ħ��������ֆ-S�|�.�D��F?�R^cc�JyK1ߘY�}�d�s,)��1N��Ų�+�w�;�������Щa�*���W]�e&}�r)"�E��z"�G���Y�v�fKΛ`���ߴ<�)��ޤʂx�������e�V�s���p(�ٺ
�K�BJ��@��쇳􄰠]�ii�#����5��/���\�=�4�"�f�Zzr���N��\��&�����9qkE�.jy���u����X�� �8ť�����Ci`�[�E���pںJ��h���k\o
���ku�<��j�:׸I;(7@����|��<��9��Q�v��J��+��N-���W�H��4�%�_k���Ma�I ?�x&���	�D�2v�m� �.��"7�	�@+��4�q���&� ���v��QM��S���4����vOքÏ����C�n-ޘl��Xi�g0�Om�Od>��d���+:i�w�]��b��L0�����>�^4��v<FXr�^ev�|��l���N�5���n�Y&��������I�G���I�U���g��Nd'L�i[�7��Bwsd�))�\�9��G`����]���ՙ��Z�X8
�L��F_|���x���AZ���qtb���Cn��x�ӆ>��N��C䫫)�ď��53$1�:!�S�����m���� ����3������Rl�h����I���w�&C͒�5��7��!H5(���phK!�u,PTJ`,��afAH[jo0hl���_}akm����3-{/�x�|�tWL�5��8^�k�ש�įWj�����M��0Z�F��B���<l�9��� ��x_@F�8ѡ�Aybn�z�lRl ��3�m*y�~(w�N����j��)ʑ�)4b��+���$�������k�s�Z�yx�y� ��jA�o��)	C���i���YL\P�L}�g{�X��x���=zM�N Bo�9lIC�Օ��3�Dy �\���
u�mӮ��6%�J��絤|�O4`�c$<��}}�T��F	)9��a��7�e	��I�����C��訩�ٍ���d�>Mz�4�|���al`�W�'�����+sYsz��<d	]j� �P�پ�a�]%"D BR��Ex��	�0nG�������ݿx,���Q�^��q3x��/X�ܵ�̒��ͳiD��O����s댘||��Sh�p10�b+jja��6W�lO.L`������8C�O���cx)�h�z5
Pu%�Cd���!`u��Oy!���4j���⊝�?��x�a�C�(����T�z�t\Tht�S�T��p��\�8��T�j'�70��D�%�
����H��v���۵�$����4�KH�&W�=B܊;���A����оQ�+���I�._��~Y5<�B,vV|C��1\�Xd!�'f4<D�G�kv'\ņE��0��@���B�G��tM+R�v"]ju�v�R��M/�� ���w�C�^*4͠Kl/�I����OU�󘩾�Gԃ,,�[�����MvZXj�:�{)�k�*.�-���<�	�14�~)��~8�9�D�8�1I���k�9A�#2r�-.SJ�D�t���"+�l�~�~�9��f�����P�՚�x�CG�h��R&Ϊh�X,��O�pi�}���b�Lƽ��q%#�����5O8i�>m��"��Q�}qXHP�s���dtWS-��'"���K�c��#�&/2~�OE��%h��#�{��ڡ*�
VZ��K��n VԷvaPz=�����u�L�k�|���M��T\��8���{9aTݿ+PJS�F3���Pd���nu��F�	�p��Rbю��$�~?�yg)�y׽�
�:��������	-�?�ϔ��<�6�~r�C�y:4G�:םT!��\`����*]�3	��&��O�e������`�ʱ���	1�T%J��IB�Z
Q!��ώPMi1���	$  ˒�>�4��
�|˲n�%��}��iB�4a�׻�&�NF�ن 8Yo�s�Y-s�]mM$1'&帉7&W,��:�*WE:���4#�H��s�?���l��Zw�2�K����j��3����Z��V�����1�[6*���S�_��-0�:�P=®8"�J�Fz6��#n��m��$��Ta��$��Ā�$��/>~��k�I���cr#��Ǜc�]h�O,rl�)BCrmh��\��v��
餕�����m/�|㗓u��{�L�������4�@���b�
~�J���yz�$4��}��P�$_�{vsJ!�=�=�,|\�f{��.D��[U����*�4+�Dld��_3��Lʭ|��)B�&!'�܍ ��ϋ��:V�W��M9�f����R�z=H)��XAYUZ	�L��lp,y@�ť(%"؍����"Y�)��oO��;[E+��B�C�4����7+��ъ�C�����~�z6��|���`}�D��1ޯ����ڪ�ɗ��iQls�UPv3BBiK� ْ��v-۽��xۓ�0]��w��#����\���ۻ'�[��nW߂ZLU͈��E�IΜؽ�&a�^�R�ݩCm�
�=h캗��f4�+�i�&��Y	�]F��1#.:Y�.��\Iz/<���粎L��j���i{�LWI��Ae�MQ�|�P����������|��u�Cv�d��%�'��c��j�]ʳ\��4�=y���nv�S��zp�7* �Uz��?�!dR�1+>r_M�ݳ39�k7�J|�h��������`.e��\@�z��r�[l�������Z����k�a�li������� C��#�˝�S��Wj/��˖�?�u�f�
�F�$����Y�]��<L�.R
 ���ם��/�V���tj���p�[�R���t�&�9-���pG)����j/��+�܅z*[��Ϙ��Ka �a��,% ׭��e;
���K��\ �m�A��i[�;�bo��`<mc�� \/x��F3%ޢ��#����Ӛ��3���f�Š(�$k��Y��_��OG�'8���D�0�a�_���ǹ?��Ն���ֿ[��gH�	�����-P�Oa�b/ �h�[�fO�/������=0��`&���SGY�+лʢ��i&gU�z�1x<��*�>a��F�G��y
���e8ZJ�^�n�@�QL*�[��
K?��f�)&�=k@�}Hϝ�#�U��ujL6��Ѥ�ͯ�7eC��dD+*o0�1�T�_��j����̳��:ٰ����:��= ��~íjV3��о!_���p��Af�A� #����X8�<�bP�R=�&��))������@j�Eb���{��/�ia��Plz�iU�_gb�95Ü��r��
����j�K�TU��FC�]�Oڨ�y�g��H+�Y8Q)9	b_fy��d�p-;R Ɍ����kGb@8,��]��<>Ige�3����T�d �DK��N��"_��ũ���r> �FC��︗�!�;���
�l�d��Yv;��)/�>VnzV���_ӊ[�io<Uq7���]���f�>S�<�S��A!�⧅`�:�޿g1�����x ��~�K��dY~�����X��΢�P2j��H��Ԭ*Ss4����tO|�rY!����Rp�$l���.�yEm󞲢񽪂$�=m��C�U��x����	mG�b�L��
�-��-�-)���bh�B��M����;��V���^�p�y�=o��W���:6��_;�����VD��|��x��O�٦l2�Pd����L�Ⱦ?e��~� ��Z�獆,W��g���3��+#7~��0��E}ϵ2igʘ�j[��{��2����|�A@C�\ ��P%ñ;������&��?���ؐ(N&�Ә�c����(s�BJ�G��ǅ�vj����Y��R�"T����˚J��iZYN?�g����.�*& Kˁ<�a�7���_�����f9(��K=���%P簮��8e╏��ŋ"��h�ff�8���Mv��<���f}%E�"���	Cm��XK#[Fل����,�<�Q�9-~�A|� �q�Ln�[�n�-D�٦^
g�&7;�X�D��L��s�5>"[C|���h��!�h�R�F���:�c����3M֦R�{=d�F�;��}I�~P=L�/�SJ|g@a��Y�
' �z�M��T��.�D�ɴ��u����,���CU�F9Ma��A!-�˅��>��� �Ώ��n��wc���;a$���CD����+�׺�u?l�l�I'2����U��k��UGP0\4�9�����>>0������n�ڊ�kl[�/��!��H'��z����"Z��B�{P�湈���ѿ�I�ø?��%���}���Y͛��m���~ǎ3��q`}�=�x�`�5��7xo�W��}_a݄�ۮA��`_����Q��`�L��*�嫵����Onu�`>Ts�?�U{h�U-V�����͔���wh���L�o��Ӯ>L@�U6(���e�ߡ3��anjRn=�~���\�`;���9�(l�T�,c�!|`���;wW-�����G���@���h����6��z��KӚ�7QDo:s�~PVxd��zp��Ud9`U+)$�)���>�	F�3�m����cH������R`%CaΞ.�ZQ�z#�֕�Vye����O"�9��gYJ��hx��BV��D�:��eRW���i�<$c3Qp��EKl:N���y�Y���
�G+��A��$ʯ�q��#g���/��_�s���P��c�E�}blD�C؉xBl��ZSغ�irj,{����tN� z���A⍖�.���|���j}b���g��LE]J��qJ߁d&Rs��!;i�����4��PC�3����t�����T���/#Fo�$*.�D�t��~�ҚO�>ny���|y�����^9�3�vS�����'<2Om���[� E���Н��z͍292�Mx�;l�8����a�D_�Eʵ�-���tW<uY�}F����\��R���8�=���z Α
��Lhպ
�^ f�)�_�e��M{j���$a������Su��g��i��>�ׯN�-Α�,sN��@I��Hڣ��=���$V�=�Eנ&�*�Ɋ&�S���bY
����|��OjԂ�v��i ���+O�p���~��VIJT,�A��y��͚���=���FJ�,x8Z��\����G6N���J�h�a������A��o4�n2f zæ��l��E�>u�g~���I5�ut�2~�H�Q��SF!Ga�h�j�6��M6PDn�c��O�[1�������nz���5wyz�
G�ow��9p���_���h�1dٶ�x�Y�߈�A����Ԣ�gCB7�5�,e&�x���qJY]�I�~�΃\�ۘ����Hv�A�v�=���RoJ*%	�����'�I�R��ͅ*�-�*�4��y�#�d�����MG�(�h8>i����d�����!��y��瑪XUL���3�p�H��~[�+Y��24�Lh@54�	i9.��{�~�ߜ|�p+��X��LV�����7�q�y�#,E��B��N`������.�_��E���9?^^Ɩc֑������9� �1
?Wʞ��ҧ��皽�'~yꙧ�>�_��N�]K�gRlj���b�FITd�Mf��"B��m�E:��=5F���wȬ|��ݍ���[>z�z+O�8~F,+7#��?p�$�|"�d�T�@Y?	����2~���/m.�fj���{�i��j!�Ö%I��t	��ʋOP��-l��o�,��D=Ow��mX˷�f)�M�U:��i�
��(�(w���Iyk�J��^�,T����B�!�[��������aJ�/�L��=�{ʣ�@�p<��8Ⱦ�����|�(��w�5���I�qB����g�ڕ�l�J_��{�*)%)��s�h�����LS�F��T��lx�o��Qe��Xr���L�x�� �����12��M����m���\Ec2�������+��aLJ����`{:�{;��	_y�W�=����e��f� �}h�d@�Wk������x���~X��+��/-(��SD8)hWK�kH<�f.(z��d�9�W��{hn@���?�R�����+~ۅh�a���Ȓ�:�|֭D4�ˤ1��e��PŁ��9���ݤ�ןL���)�S�$�!ԙn��O]��}`]
�'O[D���2��a���EN����40�����g����A��u\��"�#�.�P{����'�f����I��]D�U��fDߺd0�t�#g�sՈ �'�A�������[�#;`�nЌSf�r��?�`�? t���l�����of�F��k�Gl�r��EeoYf �Z����l�}]��1��ܥƔ��:���R� #�Yg0���I�Y�@� ����s��f�"G�����/p��Х���S�
TбC�g�,�����n����A��۹����
(������ٴ�B\�QM� ��������ĕj���oNr��n}��n�y��n���vpҮ�rC;��(�1)>����Nʅȭм�s�e 'ы�!�q̇+��F�fL����`;g���N�t6��6�Y��R.(��Gf]�h�1���A��nμu���[k|��T���_y6ˈ����2�4�����z�������C�ho�;?��!����Ҍ�_���v�i�4An��V�ȣ���;��2�h�]���m��x��}K���H1̏u��g_:����n��ψ�kT��P�A���lNf�l^���.e����_C���C_0�ה�H���/c��CNi]�I��gT�U��H�7�xdT�/� ˍ(���֢uf�w�7F�,���M9����@ U����Ac�����p���>-�9��7�{p�+��
l�ᙦ�#ǒ�JE{VzȀ�w��Nww��P���h&�L���_^Q��c��Ȱ���B7�
�Q�uQ�����'h��L�i����Αj���b%�{�-�Z"�Vu(ŉÑS���K�B�Z�,�����ܪ�w�f%`UB�5P�����^@7J��dO@،iX�q-�pR�����6��o��i]��򁀺 ���Ϊz9��~`���!ua�˪H��+P����˃!E0BڨeM�_* �!�S+X��4��l��k�w؎�+�Pk�����O7�s3���Y�=�1�Ͱ����'����@�Kި���d�;�nkM�z�A�?����x&���
Vw_<Ě�..�6����,)#�d��������C�|�%b[�G
Yk=����bTtZI�e@(��/'<�	�X�J�u�]��,Q_7���<*�h�V���[t (�y���b��U���)yi���X�=��z?e#Yj�vF��/�"��ehV2��\��ǧ��TS�yq��I�8��31��f���}�]�>�qM�9uq�qy�8b��Pt���gQ�4��ٙ�H��T�M�3��+�uN���� ǫ�dU.:��]��)�gԀ���%^u�H0w�ձ��Y$G�k�[p
����+���m��;��GُT���EL|錃��|������F��+
�ndd�]�����~�KƜHܿD��]�PtH�b٬]�9�V@�8����H��gA`A�����ɂ���1F)5yv�Y�j|�:}'��:݁Y��j���k�p��O=Kp���\��	��O2�-?v3��@u��K�GNڈ$9[1u0��4�$c�ԭ�(~�2��=�nE�Ļ(i�����YUH�
���X$��֍�#M�9�k��0ZU������9H�>�侜��e� r�e��(`o�=����P4F�i��BT��y=L�h���-��o�EX6�q�Ps�d<���\� 
����Eu����#���J�e�Ȃ�� �V���	R�Gh������(�`�rz��IT:�׺I�Wh� �;{�>b��<دC_�g�l����/Ǝ�<R�t�R�1T��Lq����������7��pJ�l[N�'�A!��CHD!�*��զ�݋��W&��|�����b���'=�O'9�'x�#��Qd|{3�H�����Z�.щ�O��G����#|*��^�u�j�Y�(�+�+�Jq��f(R��O's(qKa�PB�/�]�А�A��s�++��I+�曅\��w�ܰ��<�`���bݢkK�OgK�B��!��^��i�j<��U�[v�ߙ�����	�ߨ6�ԲA	��MA�.Q�K�8�J�ڠD�|�}�=�&j_}ca�bV��|"K���\�hf�L)�x�(������H�	f5���Ї-�B/ītrtj<BT�;�(ѓ� �%6�2��Y��1�@p�{[�e�sJ�%����} ��'�c.�F�*�(�>���y(���?�| �� >��}�btw��4}��І:Z*��81"�:�,<��/�P�d����Twߧ�*K�]i�*Y?�Nz5�X�䅝����(r��H	q��L�#��d��Z�����W�pU�'a�D��S*婷��m�����ɪ�|�Om�s�aď�a�p�h<fCb])�5+S��n�'�p���(k��&ȳ���3�i@ ��ϛ(�DD���u��|�A�t��E�u$/���.Ip�y��Vz��h��_�`�#"H7*w�:���	?[����Ʈ�-2-�{'ȴ*�E!�>�V��0�`�N��q1d�E����>V<��i���������{�F��L��ӞrXu���נ�0	Nx�s6cg����|�p?mX��ږho��� ���إ��)K����Ɇ�a�#x������緡���T��3:��cN��&(~���v�����:��2Ul4������~Mtȅ0��q��N�K01y z���'�$�'�����<��8Sͧ��N�*��7�!�����Ξ��󋩄Y�z�M�/���bn��7.��~�~�Z�H��Ї}�������o)i�a�u�waT�큠$���[F��s�Um%Vg�.����xܛ߰�F�'�OD0_
rZ�o�(1k����5�_��<�����J�Xx��,��$~����p��4��Jt���!tಚ �4��4T�5�oO�hMs�;ؗ'Xx��C�U�i�����Lz����,��M��qחA�_o�����вCX7pO�`�ĮU3��i�>L��/Ɇ=�\��Χ��3�}M�&h9�A�/@H"4,Ʃ�*�#�u7�@�&f��1="R�`�[��ٵO{���
#[��#��U�Sы8[Tr�dJt��H"֞A�;�n�
 �2� �x�?PHq ��T_�74ڢ��cvJ���/�["���/;�.�ân�6�J������
����7�O����B�����ӱ�N����=&��e�;�����ދ�8�����|lH}�j>����b��v�%���K/�}?�+�8c�Ey�����\2E�3`��D���"ͧ�1�V�k((fԳT!����'g,��`�����<��s_���-��Ӎ0�Y��%Wqt��%':�&m� ���#�w_�q���:���� �-p�o�@���Ċ�z'.��D�beԘ���̞�H5"��l#�G�ݴ�O����.�ҩe�P����C0\� p�)\z ��v���E,�a��Y�-*g�L�'X(�"r����V�[$�<DB2�!$$Gh��H��ҵEG��ie�Q6Q�@|�#D�$�ɧ���8�k-�C���
/^N03�O��,��Q�cNY-�n8+� ��.��./�"�r�HU�a���.�����#ԓ47H��v �?ˋ�?8�C�"��}�@ԫR�>�h�/��H����Pg����뙝pq6�Jc��٫p��X�9�xG�����y����{ �=�گu�������� ��-"�<��;g:��'�W�гk/�ǎcyc�UϜ�pT���o�J�4�R坰/�ET�?�^s��Q�k��g.�M��˽���7���r��E�m��qt�l��ĦO��n8g)���c�����+:b3��;�=~�36�Iʻ�ɍ���xH0��R\���I׷zg����"J�w^-�:�*g�kP�J��Z�/��9��r�m8B�[0�ӽd��衷�ɈP��u�>B=��I�F��u���Pl�d�7/ԃ(���&\Ko=U�y�5
*�B#^'�e��	ږ9�t�u4�{�q�qm�!�>�J8�z� ��ƻ��y�1:
8�t	V��O�p�g5d��m1W-ܑG�Q�RzRS�\v嘆"mE� ۊS^��KDd�H�mJ��ߢh1olM��j���51q��TX@�0�0ή�m,NL�͋�M�KI��Hﴟ2��Br�ݼ�"��{B7ƛ`�
#�_��D$��\���R	��4z����)~P�=yVʾ=G��0�11U���+C���~߼2ϒS�]�{�wc�Ŀti�{��S4X��]�}�8~D?�>�0"�w�3�L���}���L=��y���?�t\Z�!�%o6�����
�^�^��c�T?���W1���d
��FJ��h$������*Z�W����R]��:�-$��,b�9��s>��*�چ&
��gI�5q���[�4���'�_,]^���_�S2sD|M��@�f�;�5�s�{�!�.��-����s�7>��B���?C�Z1���g]w�<Udj�������N�=M�5�"{���*U�*,���:�At8����Fr3���j���2_+�I������W���NCt��#�TAL�>�S���/n�Ay�TN�B<>�５GC�^�5:XW��#�tod5�Id�U2���<�Z��+���|.�SJl�Q���v��p������Y����C~wm�q�K9�Q�E���#���XD���yL�pՌ
�.0G�Z�	��~�pt��8:�`)����)L�<�<�8���7A�U����j���F���G�8R�w# ნ��D�r�I=�GG����B<���'��8a�:s���6��e�I�V�;�#5��Va����:U�����+�"/w��f�L�����:��:�����e�2�_�����5����)i?������RS��ԭZ��5p�Ο�Z��a�3�Py��/e�ͭ*?ڏ�fC,r�oN�>�ES[9u�S`����3��kS��y4��Qv2�	�6@��VPyy�+Nפ���:�*ffN·�E����m�Ɯ�s����	Է���ݕ���8@��������QE8��Y�b�b�B����lD�Fr�	�����qR�|�@O��	�ʧ������������a���?�H�t��%ηp��B�"�m�{�����Kx���!���=���Z����og�ț��z���
2�r��D��P���>�m�Ю��\�d������Ԝ�8:�I���f�oب��-{^��Ա��ƙK�_w$^��[-R:)T��Vj^F��jC���k�	Y��_�";o����]|�5��*;�5D�ө�]����܏�ݿ3E1#		�ms�q��E@g�����.A{�	i�}��g���{i;E�Zu�}�h����~�59�oѩ_�9��|���� ����=��8��!'���s#��Oj%��2[6��#��h�]�}�����E����������w9�� �W�D��$o�(QG�R�zJL~XͲ�t�bM#��~���87���m��8��|Ǻ]��ByZh�M�����	M�8�B�� �? ��M���mи��2��M-�����┓�mE�n&H8e���Z� M9
>���w:`�/�]�6�[���wX:��mq[YO;���o��H)Qff�,�q�
M���|��pJ9�`�vM�X�L��<ږ�Yս�¯Wq��ds��1��j���,�m�U|F�u�c�<zcdO��ǽ��6 2؍��1��e�I��D�R5G����I�E�)������<�N�X�����?bi�h���(Ivsjy֋M4��� �E��`�3�V���0|>�L
�y����b��Ǆ̬rSa4��3��T�(��z�A@�l`)���/�߆�8ձ�%+�1�7�I�F8�0%����`��h���Y����ZH����&���@�=?>P�����؃����X�a�GY��%��H�	;��=�'�"���M!�ۙ�3�/6,K��1�V�@;|(��6}Hb����\�c�n��	Q}ja��r��b�L����u��$-@��Iv�R@���ܧ�C�R9i������w�}�Q
6:`���*rT��M���zB�5����W����������L��=Z<�)�{S1:(�M��ٞ��rֻ�^>�Ko�M��78�n�H׵��d��5P}{�����Jд�z��c%�=�i�~kh!�A�TP�ª��\`�Xy���$н�|�(*뽂gd5�=�u@z�s��A|pd��-%�+o�iO��1���cLk*�ժ0�QF� ������.��1*3�tVS���S�!����H(�x�4J�p�͋H:葤r�欯����ٕ,���K���^�|�k��
Aj��v����[P7B�i�g8�b��t�m|3�?�z��.sJA�{��49^'K=������,5��"�R����w*�F����0Ă�/'h�[6���RJ������}���$��FH
�N<���j���q���O.�?�&:��wYP�rs<�L�r�� ���?!ϴsσe���!��zb_.��HUj$��k{�6��1뀕�+ƈ��ӹb����$��Q�ʣ���@��pn�������v1�;-��`�%2F/�Հ�3�ҿ]� ���󾩞C��7=��"]�R��⺑�p1�9��G)���)��10ƕ`>��Q�������]\������8a`���#Z���uge��ðD�/������N	��?��xo�bp���Cι	P���������u8jEJ�o�q���c>�l�9�m9��'|@擄-�5lpi�He8sN�۷�xm����A�+���'�E���Q�P�x�O�!ї��7�1db��9�j_�%���gh;��v�~[��.��rrz�x���a��l���FpZ.�l�$�?,�t�w����qH a �MV�Z׉.�Z8�����$ZF>� e��S�>G�ֶ�� �䌙��jv|/�W0�������zj|�%)�h�#2��,��z	�VE*�T(gYZ���Ǥ�8A38 E�k@ؾ�LB���6����ncZ.UG ��@ȉ:�lW�RP�V�����pV��!TI��X��1Tg�L�?me��J�3��J�)!�+��b ��J�%a����J)-�wU���[�&��(�����biG�]	�Z��y$�Nz��j�dXE�J̮�f����;E�%*�袡�~�=��5��qa�gѩ!��ςEd�V�e�3�e�\j���F�;�$�i�"m�zwA��d�XL�-��NrOD��_���JDs��_z��苗���\�+EĒ���������Y��+fHH�hi�i��H7Yaxx�aV���"d|�8v���;Q �Jۓn��0��c�po�m�n�W@�g(ylJR�5�Bg�Ei������<��O����?o4ܶkn#��I�[Y�c�?�&^;�XnG��vM�Y;�s�I֝r���{���BeO�RHq����V�1��j/D�32.��~�(ƙ��z���ڶ��y(z�~�DX��O�y���w@*��x�C
\1�7*���p�\x��g������W�)au�Vq0t1��ʿ�\ט�Aeu?���-���6� y�kq@AE��3K`�!�Ӫ�Z�U�O�[��_��0�v6�[�ʾxQ��`W�F�.��C��`�zB��<����°��q��=��%	�n�{��0ڽ�,]���m~Fj%PE�ҟ�#FvG/����%R�㥓��m<(�#��4�`�7�٦M���L�2�T��2Dq�d�Oce���]|��ӣ�@��J��󁘩��y�IO�H�i��@!�y��a�J3����lusLJ�Fێqm�0�}+ �pƸ���*Wd�i��O�(�E^j���σ���~9!i�o+j,v9iq�.�m
X�B�[\LnN�}�"�	}A������ħk����umI��(Y�w9���" �~�厒~E�ǛbH���c�K�������L������ �����������XE�ʮ��3��-Y_�{@����%a�k��;��WR�`��gȽ��]�Ϝ�q�������hI����TۀV@v�\�=���������*�{���:QU�8�����\�HP��
��#h��3>���15$Ӯ���=k��V�k�������-����>����7r��w,�����!J{8�Z���Űh>`NV�:I�q���X^�uPz�d��*�>Vo�ڟ7��E�˓�~�uE�$i,���w�6� ��Y�(�G��c �(D�F�^d�"�%@��=.I�����M��s�����|0Ѿ����j�w�2R��L�WQGN����$�a6}jY;���?*���K��-w��o�C��ɌxVoB(e�TMܕՀ�������
ּ���Po�,f�q��v0�b�Z���/:��p�}��D ���7���+��
����f�j��ɥ���L�/�p�%�p}R��ZR!�������C)�������嫔މ�z��b�Z�x:C���
��3�C,<]� �&�����|��Q����(�$�T��A�Q*�Z��f�7��oI|����,�Ϡp���7M�=b�-_��K1�[֊O�G��\�B��c�x���[�+�@���V���v�C����`C46A ��q���['�ܬ�nT9���kY���p�q��Slg�Q,�W��J�n0p�����V��̭E���#�N�*"7*����9�kn<��ܱA������� ��h�c�f��T�R��Y��g�q�p�(G��(jaϳ�������w�U,k���cӐ46����:�+�:f ��0��L��!�y,�.p�lvx��\g%{=�{����k�9�M��7�d�ں�R���x?g�ְj%�72��Rj�à��>�W�^&���\��mgW���S���!�v�90+5���:����������tf��[�z� ~	�@(6hlO"�>� �07�^��|�~�E1��}���Hh�bq�ڄ'SI�$+�(Z<p�a.أ�������PvW��s
&��X���!Y���ϕp���Ռ �+�0�̕ #t��[�t_ۛ�r#`�ǰ�au@CNi��H��pY�"��i3�X�S�)/d̠��+���M�_?�#���������;�8~�����q��&��	���Jަ�U^\�B��g0
:;��H���/3�*&���Sl$b�~��{�!�(i-����$�$q���)��F�&͔|�3����aYnM	T����nACm%d
�w��}��m�����s(�qwN/mu��(�R�7{�s��t��S��1>�/y�-�ȝ �p�f$���C�\�0'�yT���LK�hǮL�^t��i�!{8�{\ 6�T��6W���:Pzn-+>��n��d��ߡU/ɿPxJw:��Q��ޛJ:�Yn�2����[�twQ�q�X�*�ڡ�7�!Ԁ�'�(	v�&��Ҥ.I>S��my��Q <��6��M��(;�1RE�ڹ���*�fj�U�ζ�U�F/}�����f��
z�P�H
�8i��P���`�5�t��\�j�����4<t> �R��
�k>��f*�w���F���G�'ErU�uzc���"Q��>sEʪ�
?��A�2h��8W>*纣�c���������Gd	4HEW%�ԧ�x�n�
ƍA�i�S��3¤�����$A��+Ni��	�R�4e�ªP)�L×�)֯��۶��(=P�i�?�#�!=s��3(la��w�����Rm~Jᠷ�I����-5�H;-��O��0N�~�
��\:I���!|�(���=K��n����b�x��p7�/�j�fu�(p� �9'�����Gb@RiZ���!�u�c`6�s�a�fP�}��Qc�㌔J ��w9����)[Z���6亂���L[ώ����ʎ�o�U0�W�K�a�.T	�q��/��"���sc�N�c�QB�)@�"+��"*�w�c�����ᤣC�o�fs���e<"E�o��%�����w�"�ީ��T�7f����'�(`�fC����O�?J�T�c������ʁ�'0jS�j���X'Ǒ�`�6#�&�į� �k)�qx�c�
��c�m�N��)ٱ�`x�D'�NlP!���h"��s�dD&��X���O��@�	�w������"�#���/�-(�طڎ��h4�L��zM��	$Q���Ց�7����F���#�˩�L6"�	��I>��B�u�J��x0�W� �e�U`,���<h�J$�늜T|�&A�:N�)�|������<�7c�~ߩ�J��C��~/r���
L@@g�����l1
=x�Sd/�\�A�3EpZM�`��X�y9	�HT^/L�`ʺ8� ��>K.)��G�6�6��O*4�B�����O�==���߹Vt|I���"�ʃ$1b:��&1�mq��4D�7Y�$~m�e#G��žzӿ"���_��S��n;[]�6!1��pSy R4O�eHE��v��PgY�{QW���gV�����֛�"�ˀ��yA¹{6�B$�@�.:���A�����W�X�˸`�	Zr�Kz\�W��
�C�ƪ,xE�f�����>��e=	��5r�@�ilSV ���ޢߌ����\�I 0���<�o�=v%� �EB�R�o�Uφ�\���~�4]��*Nи$���Uu�Q6�v-���"�yYB.Z��V��Fߗ��qC}��q�z�qݙ�gUG��VE��QÇ�.�6��:��N{�s�s��;�O��סl���*:+��u<�}�}Ī�}e�V��*-������=��CEA_���i:hɱ��r�[ft^NfW��#�����՟��(QX|�e��d�0������zB��v�f�8�^
�h�ؗ����uaw�XQ5�E�f�F�#9�{ԥ֞�Oz�"zN��Z�AWC
�"-a4�}}I�M�������t�o�R;��؞��9�9�+�!�����z<�k[��}an�V4>Ư!�'G�.
	�&���m�&�R���ѵ�:�g���]�GTz��_��3m���|i����ނCAdB�Z4/:�c, z�o�cB��oΦ�P�� ?��ݬrTv������(x�(�{��'0�7�Щ���� Ν��L���	J�4�.���(�=��0�Z@�7�͡���{y���u���E�c�v���&�L�� ef��2E7ʡ�9"Gu=.^� ��l�YU�l��hc�Y�'F߹��|g����	���l\�ı
��`�F႕;Rв�s&KX�&�󎏫�B�@����b=S�OU��s}�j�n�	��I��Y�����V����"Ik�$�w�w�{k�g�o�΁e� WG�5��(�%O��rez����GU�m3���՗/S��0ʗ�s"��_A���?����= �=�k9p��F:���9��F�����pő�շ�&�]9a��s�j����F϶�+p�~Ο�h�F©�~�U��r,O�:I����̵�朞��o�����-��\�e��#�h7S�yI���GqA��J>9sP$�,���w΋�/T
J����}�~�w���Je7��u.U��� �A��#�����'�1���Q�MG��nvBɷ�V�յ#��ۻK�^��?�1���M�%y�}$G����O:�{5�+��� ��V�����kӜԵ��MTiQƙ��X���-	e�Snmjز�1�W��aN)pPb=T�	��sC��]@2Ny�FG'c�h4Q��\��@8�\��=3m;�(���^Gf$QtA�2���0�P�NBݭd"�����uS4���$ޗ��JU���$��u�7�W±D2�5�)�%%�.�H�b\٦ISo������� ���������=y	.��c�&�͛ć�2 |s���L0��H���?��u[� U@޽�D/yz����������f=H����u`�'�0O�a{Xd�L	�@KA�Ϣ�J`w啃p��9V�P����錶0�eM��b
�����ב��=�=T���#�rc:�����&`hE:��|NcO�v�/��@�y����ek��tÈܐ�5d�_6����L���6n�E��pCΌ+��)0{�l��2���~��T`��+9$�� QM����p��/�-7�f�2ֹ*.��e82�*��{��X��Xfg��C��y�U�?�{B�]З]��P�m��K���.��v�X+��Q�F𠳯�b�r�����'�?X�?�H>���s�&�e�,"�����n��FO��cz�?=�t[<n��H^�ZM��Kۥ�[Vm���ZF ��3mF�W����������W芸�A.����V�t2[o ��'�xDI(=��NJ�FP9�S����;A����j�����>�|g_�QH�-�V�z�i�m�9�/��|˖��H���x����y`<F���%qH\��r�.���+m�>p�бtU&RTl�Qq�k{ 3�A���~�5��'p�A��piL���Fj�~�#�!	��z�ն��p��o�&6E��~��j���J~~"��������yv˅��3��\�EB�~
�T����Zt�b 8�-	�cv��-��tى5,�ª�ƫ��s��0�}uʍ<ͩڞF&K����Mx�:�p�x��2�>�K-��W#���P�`ƑT��,�,o-�;q=X*����z�a�V��^1w��������=(�UOg��� x�kz�1*pC��>��9��y��+_]�8j�ћ����0YO?�%��r�#�^P%Y��<V�ܨ/!x�U�x�k�s�(Q�+ց���5-�9��0;��
L�|��l]�SZ����(��l�b�������4�ֳ���v*��{�w-��Ptȧ��y&ۘ���u{r�G�	�6�2JU7�h�/���A�9J�?O���"�=�[��Q5����d���6�����$Mva_�y�^�R�!�6���0��J^�����iA�9��k
*�IbO��_�N�E}C�d�7��{!ױ���S��H��@�fЂ#�HQ�\�Gz��b�'��4x��@�o�v�܉�Qx_/�j�X�B#u\����C]��c"���.����o�ȓh�w#P�������/pC�a��ŬA��!N�	��>�ßɑRh�6� ��.�L�2��]��g'ij٘���2J�J�7����)o$y�1a������uHB�<�^T�ө�� fE��C��e�3�=ï'a��j��r�p�����ee��ہ[\�ѧ;Z�/���{��~q'��lV��T�{ツJ"Ǯw���~�x����a�稆�%v��r�Q�&�xO^:���`[N[�}�%ܚcv��#7#rd��&3����^ʤ�٤� ��R��:�-Z]o7�4w�����)����,p�����Ai��H,��9r�׫��l�
|g�I#~&6��;� ~�(�s?rZ�^�#���*�<���P�5��wjZ-Q����[�yT��ذlw:_>��T�w�^�k�ꝳ	eS���0����?��ܡu�)>����K?�I�j�Nd�L�ߣ�	�	�`�al�Bް��4�[#!�)��,�Z@:m�v����1�8�ڇ�7�ƨӯ�6L��i�|HD�i�S#+��º*���r�E�!�bE5O�0�)=1X�]�S�Ν=��WT16#R���'��мR�K�5��-T)�2���,�}���ar�+�߻��?!\�ͬl>4j��oǵB�*Byڡ �ٽc�W]�u�����
�S%)ڱ;�w;�c��]��L)���b�"�4Ԝ����ǎ������KB��M��2+O�0̥HOA0ldʹɧ�0�H�y�9	�v��eڔl��XS\fx��x��ȗ�\R��>x��c/4�Mt׭���]2Ŀ�^�
S9�@;w*�#i��љJQ"9���KZ�-ۖޱV�e��Ѩj�)��b�� ����L\I��5MnЛh�  F�g�CV�M��n� �_C��q��)����ي_f��M�d}Zx D��c�䳷��g�[%��_�Κ�N6�/����~�hr[��v�'���8�pYjx��
F�/�?�7P��i!"S�X)��J����h����+j���
�up��@$C��|�L���D$"�|�&��D�6I�D�H�7�7�ٚ�d�8��o���;��IH��mGRp��9�3�
�ǂ�6Zǟ�?�F����Eˌ-B!5R�{�	<�*��О81Ϻ�Ӝ�`C�b
0�~ؘ%���՞����#Cd�Ⱥ��� 1��4���K*� ��$�Q6C�r�1)�d`���=�D+� ��V�zROs�Q�u/t��j�9���lmJ/�<�r/�@�J�=�b�|fE�=Ӷpkmw����c�FE|�2�$�3КKD��#�D`߇HV��̒��m�~���+8�P�Gv� e�NiJkʂ�����#���Y����Il�Mf�<|��c����::)c���X{ޖ\N��n/��Zʬ������y��慠d�d��q�I2�"��'`�a��X�4pϢ���Q�����_�C��鐪5| #�uTr�W�&t�|[��.�C���ڏ����J���Hti-�0D�- �HȜ�6_�@XJ%1F;#	��V�d��)z�"�Q���QmJ"�S����i�2�� ND��Ը����wbA����a�
��������yN�\'$�id� ����ZQ����� Ɗ2���\m�\v?l>L��P���ˬ�'ws�ŉ���,�gB!�_}|�-��e�cO�ϓ����E���`'v2U ]�od۾���A��`�rʃ�-\R¾��1�{������^����k�2�7�Ӆ�L� >ƹ�$Z�e��0�4&�����v>�5�[(�"����3m*`�	>����*�T�i�UL:���6_g�@�zAU�I�|BH�$�z'O��A̞ ��C���*MQ��P��S���V�|�r}�hc_�I�1��2'���y�h�ir��A􎤾P�d��0����\�5�HW!_�D,��q��)g��r��� l��5���T9��
��Qͩ�q5J��W����=^��W�b�߂U�j'���+51�5$���@(��|_e<2�Z���C<�F�;M{�Q��zq�e+i��!� 8<�&Y�9�b�>!�NeW8�cp�<1b_g����Prt#�����;1�[fQz}�w�|�uy�������D�5����˗�j��[2���v�uj���#���꫹�cV���g���Ea_v�%������[tO%@�+����Þ>����WJ��~�/�NpUE��9�hZL��_2N�b�BJ���Γhc)]�.UAzot��DP�ѫʂ�/�k�LI8�D��Z�0yv�F�c6�����E�B�8��%��tc�7)�88�xtn�V��;Xa然K>�0�3�2��Ӕ}�������C��q����H @���v���C�$/�ս��oP��7�7�,�����)���J���$k{��r��i��:w�9,�5��n�89"u>.� ���o(���J)|���O���ws�q�)���*����8W��W�=�cY�>s��_��=֕ƺ⭥��MU�zŭw���
��p#���p?T�%����Q�8����@K>4��2�?�&��┺Q���m�b��Х>}u���"��.��0�=p�|�3J�끈[=0���9��A�Y����K<�ޥc0�+ &Z��z�u�s���(}qA_m�&󠚄���O�ƴ�"u���o8&�c�htĿ޴1����>/J�⩿4Pe5N➾��
`����H���^���0-\Ɇd�،K���g
�y���:>�'������Kl�s)��PF�eihf�9ҩ?6�%0-vw���ʊ^�Dgh�p�i��*��i����L:�ݭ��Q�vl�Y��=Qs&�g�E7������ۥ5C�%C���-G�`+���\��,��T�o/�,���K�XѨ�)����7�צ�jx���X�cܬ�Ѫ��w �)V�- ��yʱ_����r������W�o)��8��i�ʑ�.
��b��������O���^?�Ţ���0+b�ĻL�R�R$�QY�~��,�y������ (�����!0��dʟ*�_�����s�,r�Η�H�z����Kq�vQ ;�],��BȤwY�˟��Ki�#�+;w=B��)��زd\VPU�ܲ�4���ב35k���$(HԽKà�*�R;���z{��G��/�q.*{�#�ݷ�s(�n�d���-�^��ձ�����N�8^�N��ǒ���5?8+Wy~����c�nβ�g�h�E^�pߴz��nU�A�� {&6Q6u��t5�����/�ݢ��R铳0	B�n�&,��=�$c���ɺ_�.����N��[%��/�`��X����a��<�"
roѩ��hu#2n*5����ϋ���1�-���J0]�.nEB���C#<*�׽�d��ʱ ��6�|��T�Ab�@Ȝ�V�,	#����,e)\�i����Y�06���o�����0�/Y%��W��^�ú/hى�5.�=|-#xk�u�Ʀmٰ:sA���%o��C��{��C-�+>�q6���ɵs�����x4���VT��$@1������$�p[7���TGXS(�޽��r
��um}���Q��29���ƛ�o:������KȻ]�.]ƶ�������ۅ]١�L���:`��N��?�����Z��S6L��~�%k������#�6��G�Q�|��خaFo-3�˕�Q��d�B֕�}*�o��\�_��/T��������� ���C_ٔ�T���f7�-]t�=���Fv2#m��2%��l�����6���1Ժ+?v�9��S��Q�δ	�܀|�@��zdא���e'��̧w�c(��|y�M��T�&���pD��yU]�4W�\�#*�r��,�j�a"�ɏ�4��]�°���<�vxv~K��Lv�$/o����@�b�\BF�XZ��4ߪE�Y���X]=����Q�td��/u�Vl���-�^�w������[)����9MeuØ�-�!��<�	L���e[���hj�d����ΌW�C���'ބp7 4�Z��9۲�r���eHȜ�?�R�Z��,8T��R#�x=�������Pʱݑ)F��dI�*�˙���@"}O&��m(�}֏u��d�u��J����h���!�\A(�Sj���w
H���C�^��5Ŧ	Cۣ6�[~�BhY��n((b�xA��/~V��|������:�~�/�̮�%���A�ׯAB����q���9�rK=v��u�L6��i:�`*FU-��E�%�#�d���������T��'0ֳ������EYO�νP�<.�Fe�H��4��HO���ī@��7� nf	*�2>�Pygl��S��<h���/j䄩�#��7H�qd=QH|����C�M�X�����yX��<*s� K3���[�Rϫ�����Xi���X�H=vGF�[K0�&1�*�ʤzf�1�N�ջ*���mJ*�VM-�����ƌ�6w��	y��m�����DVż� BŔԖq��9E4F,�	�=�v�#)�M��(���xRB�Hz�(K�ݴe�/n�Qɪu�C�����*�lh�ǁ���.�\��
�$����Y�g�Σ��´��G�I1@��?�63����vޏ4�s��I9���+���,�2ɒ�c�����& �	ٛ0�M�Y ��*;�,���ik�Y�r�wqk����4��A&��$9g��%�l7�����V둚�!�}2�����-���*�j��w��Ӯ���F��V60���ȯ�"-s�="%�t���֑����]Ȇ�*�����Nn27T�S|'��s�!�������
�����A�L�c�/�nj�$g �Z�U��;���=�m+*��"K�պ+F���@$��!u��G=``9�9RPz���)�'-7�K��9H�"���PJoeK��
�E"ܼ��Bm�|Q�ۉ�6�Cm�ql������lq�q�xy���d'�*�8�f��A��K7pZ��c�,G�P^)���F��{�H�䪖F��'fMAcOn��=G�S0_�?Fq	� 7sT�������ߵ�Yl~�%��B� +�<�;�ϽOG���M���@�ܓ����4#Z���P�1=�"8d/��`h����cg��g�N�"��	�\�Q�
��1˘\-n׺�`q���S�Ô\�]��H��4a��?��=g�˙��q�[=$��FX�
7��������?7[c�U:�"�r��8�?C�����6(
"�UTC�c��R�Dŝ����Y���((��ΰt[-���i�d�Rr���d"���6a]Y�т�����.�Jp2K�0v� �B�?�����j���]��qm�9 !�y�&�{4����"|�v)�뛚�mz�1vC�-���"�|v��X�j�A\�}�6j�	�� �.�T>\�W�`���]�~,v��L�@(`��-\���0�TQ�䴉zyN��Ì� ���4��IS������%��pڞ�$A,T��mj�!�&(V��B
'eo=X�5T�?���2N� ��v�Kc<ܿ��vɎ�h&-=�����=��xh��p��d��Qj ��k���� /8�GnƜE��(n�m�j��@�����@F���N&�>�����o�^�Z>9E%F	7)E�Kr+;���}
�bʣ��H2@~�΄���L�FU�y���R�pA��ŏ�S/���m�kb�~ 9irz�$ū�����PLO a�VpC�x'�m�Ju\Ԗ��.�M�J����G-\�����7��%K���2{ܺ�]ZߌR0v`#!���jz�wȧvi�U�����5�4��f:D�h���닱s$�Րك�SDj-s�'ɨ�i,���_v��xY	�	nv�ATR��CRۏ Ag!�lNJlA�:�q|�K!�)��27�����*�6��0�)=�DH�K����>%;H~��rU�)y$��M?�,�6�޿y~.���p��}K�=�R��X�����KKD��c�biU���B<�OBɫ��e'�\G����h���E�����B�b_����4�[�� �L|T�q�q8����q��п�ҳ/jۥj�e�\�b�g��f�Ea�GKz�2�l�Q��i���3�K#*m�^�; T(q����IRH0�:��/�2���Xpi��F5�k��HK���?; ��^���ēt�y=)����a{��]o`��Cb����_*?M�n�	gk-x�`-��+��86��[��m`4 J�#|o�tM����
�	����s���Z���|�)�I�JT~BOl���a����,��LC+�Y����~.0y�q�=����z�_�>X�6E`��+����X�L��m��_ꅴVv�n��;*b|%��H��U�uD��� p�,	��׌��Tr>�"����Չ�d��t����^��	�PsR�9���rb
F���ix��qo�����*�l6s����
Ɛ1�y|I����ǣ��0�	B�+5�� ����+���M���7nV
u/�P��� ��������4�S�Pr!S.��-
H]}�QYr%o,����~�uђ`�8�N�s'jW��|�̉�����ٌZ��O�lM$*\�:�f�N;�joW����JN��$8�Љ>�!ŀo�ߟ�	�AO/�("C�@U�6�Ӗ��z"%��</���˃��$���f�?m@]fV��6���3;��~J���P^x"M�3���@�����P����w�f1�[V�Qv�f)IG� ɟ�rb�d��Y��!W���O�Sa���sbV������� s�?�N�G�Yj����A��� ��ʃ���}M��/|,7����Nض�B�r�sa�m�N� ��R��8ϧ��}ܚl�mĽ�N܏��W��eZ,��;���9�/l�En�۪B&�Q����dCs���ҦÏ2��T	
Ե�@�n�}��tb�-�͢	�è��g';E�x����(Bڔ��D'�z#��")�:���M���ߊq�+������$���Ee��_���iq��������Y�V^����J��4wqG! K�����&m����n2��Oj���ZQ|�	�%o�r-�<[���y�tvy��͆��9�O���7����|�����+�$z�ɕ�)B�m��Eڧ&�4k[���S��5>i�g���m����I�}�=_E�X�	�9�����ֲ`4���M ~���?��RB@� �&W��`�B	!,��H��]��D�,\�ml,@3%I���j��O �pN��?���^/|��l��}�V5T���	:�+�MEix�{�߮Ҁ+�qPQ����;��Ƒ}��Ũ��ϛ�$pD�����>�!B�^0(9���L�:HWR���c4���B�)��).3�_�P��cך ¯%I �d��������yh�ڧ�L�6}e�Q���T(��Z�F��h2c�秆n�xp��=~�X��I���G?e��K5rIM#ӂ����"7Xb��RrWZ�]l»M�H)����i}02R.sح}��Sѧ�\퐏= k�vW�v�
��7;AX��IM��U-kO��Dja�P,Jz�ol��8ue� �K!w�jI����6s�'T�e�EC���Q�>�n�o�T�5;�B@y6�8�sB*��v�7s�0���S����3Pz���5���n����3&�×�� ��G�|D�+jAފö�RU�_�G��?�@+��y����2?r�3!�X�1��t��0Jͨg婂�x���Β�l@�Z��Z�X>1���w�)�N+��^c�v��Zel5�rhfĳ�l/!rռ�N�eK��(ONF��w ����s�#`&����26u�vAJ�@�kO�r:�u���&7�-frCv�=%�к���r����5�w�L:��?����^��jHkDF���O����|�|����x��LO4����v���Y�aI�,5E���E���T8GdG�p��^�	����o?��#���\�a2�u+ܑ��4��g�����ܮ����,WEώf���D�`���Mݏ�3[�n)j]�j��+���a���j�dn��τv*Nz�w����j��>�C�.��52�c��?�Ŗ|dΩy�����j���N*��}��SX�ÝΝ'Z�y�'�ea����j~b
b�I\�9�:A�媣�;���VP�$�C��K;݉TET�Z���1ltVy�`��wlM�]��l���4*6���v�u�Z֘3���;&�1+�q�%pK�8D-͛[p��b���yU��y���i1�o���[�-�-�5|��,>R�	$;&N��\5�M�� 3g�01~
�M�M��Tdl&v��Y�	��n��f�Inb���!�0�N^���_�Ԗ^'PxA�T��a�2�,�Bcc�����y��`_"\�t*�5�2CU�a7�e(te׈��ι"b�3� ;²�-/�vBӥч��Τ�d��W���\~�L"�5�L�a����.�.���~�2Qѩs����* vD����$S�>O�+���^��h����h��fZ�^��w{�l6l��!��͞��^H�pڔމC�f����R@l^\�t��섏��"qjj�R��.���B]�8�7��>p��)����t������7׈��7T��#��ᅣM]�l�DaIQ-����*��'7�EvRT��w16�T����)
�:;�Gb��s�7Q<1+�5Ou���U�ңBwǼ��0w�Iu�d�M�6k�87��2ԇ�+vYuT�" ,:���$�B��M��(����V��z�߮����K��5�rQM�=y�bh#�X$�'#���)'�&q0 X�XX�KΠ*⎥kB#!'��=kx���P�SZ^]��|�ը!X�yl�`5~�t���(���ׯ�8q
��܏<�]�[���9�Y��&�A|%��&S�.����^��]RP1'�86x���T"Hsw����Pk�Y�t�=M�'��ܟ�w�D��Y|^e�U�mYg�{9(����,`.��T �-��An�6.����j(�t�C���/�U�NzM����P�>���uS�*�m:�+�z�߿�R��0��8"�Y��+G��Ƕt+ZI�҂|�.���uh�<��u�4J�pEd�'v�۽Ӫ4�L]Q��1MS~�HtWZ�H��|�[J�qhu��.yO��4���a�kΛDK���H��X���3IMRO`�@��YQW��`]B�S{.� =ܐ��"�(��`5%��:�z� �T�����E�i벴�"z�z�y)ၠ��Ƚ���l��ݷ/�U��2Y�Y����6>H@n��\�^Ρ���`Aݓ������-cl���]I����79T�Ǝ��[9V \��z�ye�)�pn{�`�	�1�(eG���y�d��.�Bz85�%� l����D�J}��M���^��ج2 �f���zd��\S��Z�����jb�D[��vvs���Z��g���"��E?�+j���@��(獍fê27뤪��Ro�����H��]�¤��̶�\Ԩ����jݩG�h������?5�6���\S��JK}��-�/i�{�{:��t|��G�|-��p2yT?	v<`-ƶAy����p��l�~5���4݅bo�gX�$�Ȣ��'S*�5�̌6�v�^���meP���2N�f�~N�<��OB���j�^qB���Ŵ��@x��a�A��PW�vAC���ȏ���l&uY?Ѽ>��ꅤ�ϊn���C'�4�ު���#�7���&,�QA�O���Z✖/���h)��
�N�����?��$`'�MO	Ά^X���L?r�O��)6=�%/�c,�ۗ6�-0�`,��+�~��"@F��|.���1m�����>̊DH/�s��ZUE�C#��@���������K:��zz\���噘�����]���:�9�,�+��Y����8+���$�����S��9�I=c���u�yU���rn���"���6~��Q��2�%��Bp[h{}�rUz|��Y>�Y���T���0X����[�)���Ӌ�k��<�E�5;�����[ޟ:�Eo�
p_%]�~�l�ͱ;g�#�^�J9�Ɂnm�C���K8p���~bC�bʬe;k���
�zI�W���=@�1K��/��!��5��y]�/����GN��b;��ݵo��Y�kО�Dڮ��6�&����������M�aߙ��-Y�"���؄��O����{b1������V�v���3�f�ΠZ�IS-�5>�|�O\ϟO��kM��e\�/��`N�Z!��ˊ'�����ڍ����U:��"�x�=V�Y_���Q�%q�.u������n0�&�n+v�lt �!��7.����<\�5����{�O��ș���Z�2�s�o��MK���mv��+�	���Ũ��X�"�k��4�7O}����r�k���-{?��H��ŝ���۝�����0�����/�T=ĘxF�B9��,�:j�� �$@.y�a2��o)��o�k�� �Y���^|�^r/7 ��`8ˍ��s�;���Xp��:���� �֜2��J/܊!�"a�����BJ0�E�|n�ڼ���w��Tbs����&���Q/��fI&�Q(@Y�K:����RN��5*��lS�L�UC *�+�r� ���)��^,qBx5�3����o�Kw-�E�5�:��F��{��֒?/�^����5�5p�i�t���^�?X]�%���dN0YRؤ��$��07�E�^����zq�����I<u���}�å�����FH�&��������N���h7�
���O.�`�Qz"�s��f4�� �z�%\���v`D����ӋZ~��7ڠ�cm]NE��Rb"���$M�AL�r���ig6\�@���[cj?_���:��AI�B7��0Y����m����^5؄�����I���Rz�W�j�#1�Z_;Z f$dVܼ?N�w�A�e\���7�lP`��l��V�y�b�ϳ�#�-*���f�)-��%C�r|i^��OF�IŎ�����	m�>yO�>t���u���/0��g�`�0R��1�*�i�}RK���D���^:QTD��?Q{�0���T�x�6ҝ}���{w�\i��j��c|�]C�$

�D��:cr�a|�gt!M5p|��p\,M�d�����}I_���P˙�/�$���֊#1_E�KkDoTkGk&k���TJI�*�-1#��,����=�X��r�-�4φ�G��m���,+nw�>�)JI���Z=h�h���$�߲!Kq��5F�/�%��~h�������bR��vIz�p5N �´:�v��Nf��I_R'���r</<���CV����CW�aT���%�c�(�/�����jl�5n���������Қ+̢�!���uk��P49o�rw�b,�K�2��
��8&[h*��)kÇ����=S�Z����x{u����r��{k�y�1a���=r��#�F4W7��p�N�-d�*1����d\j���^GQ����^y߄%��y>���~p�J��yٖD�Yi� �³�΃�Z�L
�￘���zrp�GƬ3F��D�Y���	�=Σ��QH��أ�^�v.���]��$�C���"J��ۊ�����5u�:��M�[��}�O�43�d-���2�>g��H@<N4�V��|d�/����եr�_��8�ŠT�p��n�2�|��"������0����E��I�"v.�ʋ�N�a"ʞ\�pX��|����d|�J�&ŗ�ݮ�����(�1����:�`(~�����_ٸ��
c
ۈFF�4=���_��Hv��`�!�Î���p�^�M�"��tm��hHM�d�Snj���-��u�E�B�A�#��
V��.ΡXZee�;��(���=�z��p�Jȓ����WL�{*{WI�5|�L�!Q�:k��T	2�g���u�h�t�IV�f4g�����m��
���-d}]+*�F|�7V�3-5�d~~���R*�)QP�&1��C�@2�Z3Ȣ�#�N���)��-%���zgZ*���+��;������SOo;�o�D��%I���tahe�U))ô�#�����Uz��{�w���J��x`�&mZ�c`�
p^��_x~�0��X���u�=]�ML�a�\���U!�La��lŃ{����:�j�ne�#�K&�7��;�HԂt�Oz�V�k��Х	r*�XL�t��C"�$�<��d=#
p��v�[͙Ub�-�B��7���F�ﱍ�]���%XwT��٭Rw�S�1���|%�
��@�
���,A��ɗ�q�@Q�(�Y���*�y�k���Ȍ��|4�X��pW�8a׆�ɓ�K�h��J&(&^0�AVTBzsG���X�⹓ʅ���������v�~���|!	+i)���u����o�S���7ڃ`t3�b8��l�]⃯�K���9�h��(��أ��4,��
��j���#��<�rE3����sdFWR�*��b��{s�9dǿ:W�&Ǯ�> ��إ���r�7�I�R�"icb�<l��ڝ�ư.7���O�@ Щ�'��tT��8��yˌ/��Lp\l����5N�6$��J�1ڗQ��[�4@Cc�#�|v?e��\.v�{؇�d	;7�����jt��2yg�p4���#���H;r�b���0z�������J�\6�j>�B���R��S�X�a�8��u�(�`Ro8}��DM+����{W؃�b�H�ˡ�4 ךуp�7�}�
*�Z2��.L�l���5p�N ���J�֠�f�Xh�g�
QQ��	��F�yf9�A�]�ȗy��<�Â�T�|$�w:�J�;�m6f��l%�~�Ta��^$��b0w���f��1����	VNV�L4���x5!^�$���j�U`��cAj�(�ؾ�̔l�O΍��$�x�c�<GH|�`�s��ux�i^�ε�����a�ȉc��Q|cV#�Vb�d�f����x�lK�g0$�	ED���t\]��>�g��_��"g�Ƕ1?^����K0Ikk�
hR�b�<,>g~����;k�sl��؇��h:
�W��G��f	<�X��Q՟���Q�u�L ����T�;miVj۔�����2��Jm��A2k�vR��d���W�����N��f�Ѝ�6x�7J/
\>Kx*��Q�� �ނ��d��D��SbF��ۜ��t�Fв^.N -�� �R���^x^��`��\�{�p 7O��N�n��W�*�����Z#�/�C5�y����[��_7;����̀'�-��Y���!��&=�M��b�?�ն�¹�*�N芼�\�3e���	,+'�q��LK�X��*�驧bY��%>���s��6�B:��OdRy}p��<����ȶt�!X��a9�����ޤ&1��r"��(��)%��v^�q Ɔ?w(�K�./�xQ*%�&�����X)F��5���{�3�����?�F�8@���$�p=/V�LWΕ�z�)�f�d�+�����~'�RjU��犎y��>tÿ��|�'��]����?��P$Pԓ�i���(MkX�4ee}u{���c;T��*�F�WL�ʉ|��V���j�?�������"�そ���2ݜU�w�hs������B�Z�Rr�_��'��q37�!A�W��S�oQa��4�4�$�<��&�����u��F���Hs����s&�j�p4�dD������}� Y��f�-��شf�{��c��5X��w�����=f�2Ԧ��E��jQ�P�}�S�c>o��O�R�aFK�|��~Y��2��J"�E��4����>ڇ�0a��g�:7��@Z�q��$���}��� �*�S,s�|>�f�I���(Bo@\U˓�	�[�e��V�l��h�^ԃA��鏺��~"� ƋO{Ĭ�R�����R��G��4�i���D?,t.�}�ބ�� -������iS0�^Nɠ���<M��148�wr��s�grf�Զ��)��d"�Z�A���&�~��XE�/N|�]�4TY6�m�q�݉N�UܑOyE� 
�
P�Z��wx�)�LG���壺�G���N�m���0��@�g�%͈�f��$����~{*��զQ�U�/$�����'/[K���`�țH��N��UC�D�b��i� J��*I�;��10��X�dr�����q�ʁ-s�,=Fԁ4���<f}���&�NN[�+M���9Of	s�Wk�{.dpb[;Ƒ�LLⳄ������*���q�[K�V
íjWs䞐qW�P����e�Mj3^E�L���O� �p�۟��8	��FK��<��zk�0��P�����N�1J;k�Sr7������<}��vs]	A��)!!���t��u���v_]�n'!j���u�EGS�4�^��%Np�e$}���h�n��B�i��i��BX_������x�J�(!B�<	$網�%Ք%�4��5`� ��1�� w��f2CkA�{6.H̢�[H.�Nl�}@�JC��;
BR{�~(D�C��{LYx�s�,c���x�F��K��;��	!p��8����j����n�*�Ϗ'{�Đ��L�\��j�U��\r�vJ+3.J�������s��j|!wi:���v�����7����ͯ�s�G����T.��F�ǘ���G�[:�p�("ߩR0��0���D�u�TW/5WI�
����CW�&���ռG��Y�][�yO�~�p�"` ��N �l �f�\6�+++�+�0Қ�+J�����"�E��b8P�$U����h� x@&oSL 1���U�qɤ_c5���.�� Ɠ"/�����	��qMA$��`����Y�p-��|���[td6M�QS�b�����^ֈz`�[���'���#%я��M ��t�- 3����ۡ���뿒�=�$]�li�!�Ox�(�F�r���z�i]B������s�DB���q*&�:���	qb�9Q��B�7'�[?<'_,��h6ymn�t4��e��KQé�<Wr�ׇf���d���eY���:ǗT���9I_�ɡ�!�;�,u�E�9�v��K�����i~�4	r���ٛ��s����Sz K��a�t��)�^��@�4$v��r����+t:�7�"yq���*$�RE����:K�Z�]�Q���nP����,����d�A��v)��a<7=Vl��Y�s��OG��6�|�_L��]�,i�����e�
����+��UZX]k�P^���ZyF\�l2/S�v.�
�%��`8e<s#�R�qYxR{��}��~����ï5�����ƴz��N����~�GeM��kxq���@��v�[���l�������B��Df��%�r��w35�Rxa6�G̪��m�MDI�o�{롣lg��7�a�-�0�ai�k����	;�7։߉2��>5�͚�Fw�?L{�U�F٘'�7�N�щ�k���#���B&"��;w�?ݎ�`�� F�n�J�/�ʒ޴��z�VFLW�:Սw{��7x��Ia�]4��gfb��4�a�B��n7��0����</�a��T�y�d�G�d��ѕwl	��1&[���>�������dLH�̴����١��E3�KQ"���_��.���$���\�3ft�+}8��@j��H
� ��h�e+��e񰋁�ArL�}�Ͳ��lv�-�����n��\��M��z9q����3�H˘P@����	���� �&\,�0Yn4l�;��4�o���-��z�Ē0K?����p��
|�nQ������p�CQ��A��� \ �(?�@�d4���ӞL�����"�{��^ش���f�����d���%��ꯞ�߰��u9�WN�}Й1���{�`�3D9Yd�\��3�J�H���N'����Q�F	�hE��ұ�YҺV	U�c���ʝ>��xqSO���H�@6u�л�����xa�; �չ�Iz��������g���tIz���:�V��b"��<{���r1@k<�9��*�̫2��s���vĖ��bH^���"x^Ee�W�|��,�n��e�K<�Xk@	���E~"T������ت�ZB���ɝ��m �bpx3�TX!kR�L�EQ�5�9쯷; �ڹ��))�L1�	c��-���<���(���vw���i�,{��qߩ��H�7�1}���M��U�|#�b�A��xֿ��զ�5 !��Ν[DzIl�bXNG�7S2�.�P�:�q){�F*1교f4a[
ʍ�m6�us�KTpۣM<K�ʃ
'�g�E�wY��O
�aC��f+�o0H����[�O��K � �T�m�� v�T�����Zk
�}a�	c��*����xfg3P_���f�s"�&��W���L�!ՂT_�~����j�o�=�£�z�6ϧc��}/q������i:�nq#��n5�>�J�x/�[3?������#��W�s8~��M9���hl����2�en�wOAY�L�O���2�y�{p"+��%�O� �`s�q5�����W�ͫO_�l0eR���qc�C$8d�l���}:��Q�Z�)��ܷI�y��Y�S$��c���U�,}_'?A����s�������;
rቌ���K&U��[�[Ǳ2: ��❗��~f�l{W�/7.)��E���vA���FL����9m	2����?�.G*_.�`�9��[�6o(�����<�X�]x�U9龜dB(�>r{wn�p��aOj���M� h�F��m̴R��O�ք2���hü�iN;H��"_��NS�������tR�����L�`iwۊ��?��,?C]�K�aq�ّ��B�ǻ�����s�&��:-饙�>ksB�/�{ +H�>ӭc��rT�퓅�R��#0�-�0?��.n�L�H߾O�kTH۩(��ѓ�����9�Q{gS��<&�!��m^�1��d��ɰ��w��Yl�g߈f|h�e�x��/���Dh"ph(t�M���s3p�N���O����N� bR­ծ������o=���J;]���É��/{e�����w�����a�[�A[�5��%�� "�@�6��U��`k�)�D����xi�������/�I��r��/���Õ�s_MZ�m"���f�k�?��\ܗ`���U��*�< �{W�'aۗF,9�f����ݷ=Ϳ8�$yޓ���{��fA�,{R+���G�é�ߪouF��G�+U�H��Q���f�� :�J�!��(��8���LW�����@��^0r[�L���Bo�b�/�"��0��o�!w\5%����CAOd���sa��G |U�)=7TՔ����"�_��W��o`�@[�<bզ`�3�i>��.��i��L��%ɪ%rSa �A��[���+�7d�Y*�";�pۙ|��<��y޼W横D���)�R�5�_xfTa@U|	��y�@��KU9�.%r��O�4G2��F'.�OQ�ӏػ�>�go(���ۯf�C�~,*��/;&����E�ANt�в����������B|c�z��~܈~Y���WT����h����w�q��/0嚧�_�� �l ���p��q��
V���d���������FyO�YX�W�-�� �wk���ܸ��p�����+.]��y�V��+Ƹ�P/����)��q|^��l*mM;����i2��O���Y_n���0$�sa���ʗ�\)��1P%{M�O�/�w��;A"W?�&7�7����4�kh�T�0�T��J#m�&���g�)�A
_f�{±���B��F-u�)�$wȚ ��\�sd�&~� L'�˅F[#K��~��$��0�� ?�'>:��6bǑ��k�0T��D��[���P/�7�xa ox�T}�����!��$!�	���\��2|d��s������ya�Xw���=�_iT､�2O�<Ι�Ö�(+.�.�]w�� �mS�N���4�_i�Oe�4!'�� �����i�Z~�\U���它�fjI/�1����ˊ
�u���Yr�+�Kr��hb<$�5��ÖS��r(�oo;�.���t�|HP���b<�P��k87g8XMAI\����_�k���h��\���h�=*J�'�q�Ba���n��HW��,bze�F��,�����J�� ��qm�|hp�����#iD��*9�+��C�TX���@��u��W+�ݗ�����2��Yu0..-����ZQ��z��	
�}�j[��y"�������SK$H'y�d-9<���*�yV\��0��f@�� ���հ��@S#�Π�g�7^�p�����GG����U�1��k���d��@K}5(�+2%��K>��KD�G4D�&�9����^(�u(���E�dU���/ě8��iĦ�"ǹ+�D��o-ɫ�����t�@-�o�������
.� H]���sl�G!���	vZ����$EF;�N�q .8�N�[/+�+N�����B�bI���X�5l�<�g.���A\a]�%j�I�`.}#��R���ɕH}e�@�0��C����@G�Nג5�F9��Sl��3�qi�n�*
�,�����3�)�t(e�C�.�j_�>��p9���՗��@����_���X�Eg0�V^�$G��*�3� �My��i�4��i�N!歽"�i�d9�v�}UQߞ`Fס~���^J�(*4�F�I���G��2�z�q������ؓ�U�o/�}�W��J��� h��lx���9B^��rbhD����jH3�Hq������J�tL�+���	�F��p�P��5!�=�m]�t\Dl�[� NK�;�Oh��\��l{ 5#+Sd*v����p���JRtԐ%�p���N1���G����H�:M�̿��� �_5��v5~+1N�t0�q���o^�N�4x�V�Ĝ�+O�3̌a�T�#L�E�8��|)�9�q�Tf�2}����B�ɥ������l�oOsX�V{�|���$7a^hUKN���:�V@��E�6�����
��Y����� �����Y��Mnrm�}��=3��k�=�>�<sQc{O��Zh��9�!��q��@�[GZz&�ʍE�	;�6����CݚX���ω�Xcm���yF'�Z��{8G�ɤ����k
=�bu��sҢ�!�k)��@�.��Uꆇ1�c3m<�����E:n����+Wt�F_lQJE�r�/�j���u�$G�Ĩ�"bf��$���&a◱q#Y8�ꮯ�;��T����	�M�bG����j�OG��"��'�����t+��'4�Kn�UZjHI����ͯ�[����j	���֚�p��o��WP5;r~���;�1�_��Ӆ�a���x���?��k�s��� �e�����V�M�/���Q�=���w��5��:�y���T˨R\f1q�K��������s�7L���Ԓ��Y�p h��b���u�E^���XPhyu�߆�����4��yZ�)y2��({&k�c�Ԫ�.��A�Qx
1�d`��HMO�I;��LW�X�8���U�&!ND�Y�����ӌp�C��3
�YҰ���wa,Z�%�ʊeӟe�:c��l��c��k_.��:�xH�R�����ۿ Vn�6��`��M�b�.��j1�=����Z��,l��T����bk�h��g���<l@�b}��"ۆe�~���ww����N#����/�4�?:��>z��趻��ΝL��T��q���U��S�jv�Rc�X�0J���ț@%�*�yLю2S�:%�l\=�L���V]�o�!�s��"��W���]���������-z��_�誵ڒ���S��?>������T/-휬(@������i�	(�ogwR�h�eڌ5��fmJm�>�|V����ڰk�`��ut���l��`r�������c؞�XJ��ò��T���6�Ԁ��)�.o����"��7$�9[R������1,� �2��\��y���4~:�
éҋ�3�C��s2��ٚ���4����m����7�?î���4`�=QE�����ՠ�O}�S����s�<ZD� �����E�PK�c�����|hv�}~F�f���3�=��j҆dw/R3�6<�P���A��iH���5�H��$aC*�ߌ��-��ݘ���EW?�d���	j8֦�&�!���)',^]HX���C��3����R��M<YTJ�{Bt���j�1�*�c��̘VU��zyĥ��N��U0)5&���g�烗�S�~�OZ��O��pgc���u��U��*m��G�Zq�"���U��r�(�����9)\G{S��]�vKy���_�\f$G0P*��uq	�0�&? �����x�O^6^]�`�K�Yșͦ��|��K/M���.���1��n��#@��/Q}!��A���^��F4�]�4אz�����0Yl$�A%K�gaCO�FSCCt�>ǎ3�^ߐy�1�M�{ms��-GXw���`1��Y���u襹����ҧ�����v���	ߙ"�ª1,��l�^�N�դ�-��a-�����&����u��q�!m�yx_�z̠����Ns�Ga�G��(f	cs�f�q-6&���m@WS���F2TmB���Zk�7ҳD��CDJ�������0<�O��t����C���qY�#�]M��o��|�N+��!g9G�wДṢ��L[KD�'������X����,7�P�Kg�|iv� �Ѥ=�r�2�1�|;�C��|�V��lD�4|�Ey8�Sϲ�E�P�٥�����6��w�1c���>>�j���?Ut���)�}f{c:�6M�5�r8�^Ae /
�7e&:�Wp�Da�&�����Y,L�5��SX}�g��^�L(<�eQ���j��xY�1&�*��r�]�;h�Ɠ�#CJJ�o#NHT�<K��J,��l��g}���i�Ä/�r������ʐ��P�t�!(f&��(: +&`��ɶ��JFػzK��-x����O,��֨�D!p/���k�A�[(�.E��
H��V���d���)�G;�5�Ç�*"��
�b�&_�Jp���x>y*�:hSE���}b3	�m��{o�2s�Js��,	�V$�B��	�7�{1R�=q�����D4�su]d�ND��y"wz�(@�ͳ҅�ϰ�F�wO֦���i��B�x8���C#���r�E�������B�br ��9�c��B4{�о��Xʘ�51���,�Ě�p�?�<�=�g��7K�>t�|��s�K�	`� ���	��95���!ޥ�&�w�.�)�K ��V��]��=�Jq�x�I0+�k`��8[�ŭ"Py�ko�wZ mKo�U�!fԠh��7����f�T�����\���R�H�L ���Z�0]���+Q�I��E`�(!Ϙ��?L#� ����V�����ڊ��qO��q��f��y�� ���r��:]���εU��{f_�r��@�Q��ڏ��J�Z��v~2O���)�cQ��)t�Jj�]�͍
�IO(p��歙�����v�"�O*���{�Y}Q���3��))Dw��r��_t��������Vx�#f�\�\Ɩ�a\�g�p���4�_+�]���d�Z���" ����ڎ�E�����t�D���eo�r�i/��@��Yc�j�ä���:جRG0�U��[�v��ʁ�{}�J�Ƚ���:>=hF���~d�U:D�ĢQZ�Q|��E��i��쇁;�Y�:*�`ޢ�E=�7י}��f�sm��֠�P��+�Iv@j�D(��h?Dc�nГ�~��C��Go�+�%�����q�������MJ-g�����0����V�A
j�ޘ'���ҝ-���u=ZV��e��={��L���d��=B����v9��8jQa��V��a��h4�L��N���f�CB������>篨	J.�H�s5����JJuӛ�ﹿC�����2�I�Y��^����ge`?�Cd�*$;�N�?<`:PeC�~ֹw��@�}LiL�n��#Z�fR�o�������3�0���V�\N��;ǱV��r�M�V�/j%W��Ǭ �M�agm'�WK0����}{��!/���,P�',��ô0�w^%�k��V�^C��7�� �}�{�%��ˤt�o�򮢤�--��HG��)m<���Zb��i�� =��̝ફ`����&��X�F��!�w��M;�8����;۫���X�Ś�X%��:���0�o�H�r�1tCK@᦯l-��� �.��๺��i��)&*��W��J�����;d�RZ}�����"P����>��"�q@~T���x@=ԥ�Ī&[����ҡx�_�Y����њ#.�&�L�yTs�f�������D96X`2$5�=˖T�h*7p@rZS'1���Lk����~���Y=17i�n���7$��s��(Jc����i��kP�/��W�<�}.u鯠���W�,��=i].�Ân�*�i:E�<�$�M��m>�,��7�-�Bݺ�RHP�Xq�~G2bO��`��-�ˣ��2վ��q��
׺q�N�U;Qbl�h7�c�����ؗh�e.�X���L���F���£����T�������N�=mwai��@�@��ۓ?G�&��O�_\�6�j6d�ɹ��A���ׂ�5���FP��5|;@^av�22"5���ϘQ6.J�8X��e�v������
.��9M�4�\zw�˙���ʨ.�Z�RC��֘�v��>��pH�ݍ��܌��IhG����Ł<P;�7�e���L��2>���u9|Q�|t�;5�ߦ�Ϟ��:�U����=����C����dd�WO=u�^�	`��:ҝ�c�����9���֕ȿ�{C���|�������-]c�da�'�ѵD�x��t��@�rC�Z��� Q�2�@0PϞ���� ����X� H���Ӌa-��:�f����uW˭��Fn-kx�z*Um���a�|nu	,@ZW�޿!��)T~�͏�x'��D�r���G=���ݱc���q�p��P�b�l8�C4��`��7�9�)J(�����&��	2H�O����h9�$��0������0b ~`���	 ��v�ވ���<�%�z��Bk��F�],��d���1v�\f�;H]���X�.�J!�8���b�S�.�h��t�o7ȧ7��Is<{�;�1t|)oS�dW$jhu̦zĉإy?D�� !W�+�����smӏ�{4��\�
���.}����=��/�n��d�#����aEq�vB:�)j���`]nӍ��p�cK�f�����A��PV��G�M�7��#.msQ��!���t��ۥY^j}E@BeqK�K��_�]���3��x�,u��ᖢ���4%''ò�
(U
���%�5�Y������� 5L�H���eZ�����"�BVOX5�*W���)xխݣ�����e�q�%*x���Cl�����T�'|�X+�ں4��{�n��bId0��ɒ�?2�-!-ST�W?d��@X��6K6I���@�,��:6[�˅�|7�&moh]S+�G.%�_�]��/�S��d.�ɮ$��Ԉ����������j�G-B��d�Bq�����S�u/�"�à��G��`�Ô(a/̈)�1A��G����'44��E�i��9P�F�;�k*w�k��D�Q�6e`u]���l�z�98e��U�
�q?Jl�%	M����H�����UT�A�G�ڜ�nC�.#b��I@��7)goU2i"�Kk}���nU�ZŔ3�)��:k�OK�8�Re��
�%�6ڬ���n���1x�����ä���0�v��-d3���������<���'{�x~�,�˞�\���A#uu'G^E&Pik��� �kc�q�����I�y��Y�ة���U��>�u;$��-a�� �r3����b��+�劰N��n�9���A��̦bX�g�K�xi�"��/o� [-Oz�-p@��2�M�4��p4|ƴ�]��G2@,b�O~�N�͑�6�M��.��5O��^������"�[^~z�/n���w3�/.����eR7�����/~V��_�����I�;ؕB�~Sә���!���>�B�(�뱩kQ���5��\��uF�gF)�(��phJ�^Ղ��u�=�	�b��p����쳭� �`�MЍ�m#.�պ��iu���D�� QF �!p����d�?�l����Ŏ|�9l�f�a���M�C������!�\�L0V%^�pW�ΐ���
&���r6���Z���Q���8�I4��uw!�L+�F��Uң4�Oq/�-�B%HҲ�0S�m	B(�4�4�RՔ���OV�A��7�!j���W�GQ��j9%W��	8;}�)GQ<4_�0��]K]�Wm0֋�۾�.�@w/K����gI�f0/A���G���R��MI��	�"�lƃ�̑�S���+�*Ŏ�%�5�}7���vD¦r��£�(T*$�I���.:��C��h�Kl=<|��%t�(���))����������!��O�rK�.�P8���KH�fwrqN��~�5�`�d�����e�Q(Y�;�TK��%�����W�n|Tpip,N]r\Fmj!2�ϼ�8�c2_U^M
��d�����.�'�S���+�䎊$�0D��d�j�<�-)Ry�
q;����%��.XH�DȒ�ᨐߗ �xt��<��ݚ��pб(�z< A�~<G!~ab���#	���L:.��X�\�z!A�)��˻�.��zZ��s[���&�'n�O��}�ɡL(��T�*6�x5�0�C�14o���Pb����`ODPM�1[J���FZ�?�#%�h�|.��&�����p���_kJ�Ք���"P�����靿tl=�ܨ�Zc�?y����zSp�m�lq�(�~��I/������ȼ�|�kI�ߘm�T�5����͗�,0L`�>�3��nRb���֙hO?��ZN�;&H�X�_���	��7Ȱɞ���ʎsZ@��
G�e���5���$j�wv�W8�9�˛-�'$i���G������(���� C(>/�A���M��q�b�!? $tD$��Ih`O��x�t�A���$��Sd�ٻ�������#�����C�2+l8�X"rǴ�}m��J*M�`|�$�"̞�	@00[K��a�H_` �JMx|��Vc��G[N`@���)��؈2���� k?Rh	 �DСk*��T`��;��Abd���TE�w���&�<�S�;N�»E�����dpZn��ޒ��1�]ڎR��a���>	�o/Q��=���䨏x���3IP���6ui*6 +$�dS%G�3�	^�~c�MXՈ�}���5\�ȁo��R[��y�9����Oz�ę�4�Ȥ���e6#����^Ե6����������dE�[����~^���
j�~�ĬX�s�H��Z�UI��t�=rWp8\)��Y�63U�6%"�GsO���u��J����rW��/utO R^d?7M;�\'�\�8n���K�`������"���a�V���(�A5m��%����5����{�[㊀_19��i�9�hZ�y�7NS|Z��/�wR��<X�L��8�� �=�[_i�}���uaD]5z�>���P�9��~yߝr�[� ������@��됥�f@o�pK\.\<���|�sB��噐y;�%��� U����˰�h�@50��z�CT�!�36F�HS���=���8��a�<6������G�f��V|3�H�@4Z�J��!~���iN?P$i��X�h�q��8�_Y��*�X�F
�j)������gy��p�B!�T�HХ�yu�5���#����Rp�m�A�&����A�C�>+�P����^�nT; ��Kf���z���4���,D|U
!�rd��f�`�X�݁e����6����Z�	�������T�#$)'��Ǒ��w�i�Y�ʺ��H��Tk^�����J�D��#s��M�x���� ����d:`<�'�
����av�)�g��:w����[	8J�hG��ą�CAL`BUۥIsŞ���R�}����7K�+~��C�0�$G�W��U�����i}j�xm��Y�V��-VAů9л� q�f�����~fQc< �
��J��RHF)�4O�Fq���@�{׽��(=��ǟ�J��-9��Ql�j������v����gQTLH���R~��:�ld��琤�HE�EO�=Zn<:�W���/�}�<|���w��^��s�s�����w&᱙=�k�A�cYacP�9�p?ѫFROF��@>�b�~2�n�� ��`8�~G�kH��%�>-�8^��$�����RM}܆�
��|';�YXφ�	��j�W�<�c3\����}�J���(�|cw��;e�y�6��:���?s���L�L�yB�"Y�۱�k[A�z��qg��-e���!㒯��~� }�e���d���K���6�<N���B?Qjn�̂�K�����ZV��?���?�"��Zcx��d�;�|)�kߜ��1#��}���n(2L�+��;}��(�`[-:�<h�l?���(��D��W�g4���	��%i?�lP�QD�Q�3O���j1\������\����GǪwHp�=m���sc�3rfgx�U9�}tܖa�i�u-(���^Bg6P�պI�h��-��Ev�J@H��E��a ت���v*�.F���Ff�\�F;��c���ˁ(	�Eev����^���|p�B3~��M%_�����e���a�B6��k褉JC\�5dG�M�n��M�I6-�sD��}��C�Ҵ� әhY( �U��y̰W�9��R��˵ �/��'�Z���)(��t�f�i ��rÑ�Ҥ�=��z)`��pC'մ�ׅV��s����:���-��_��착�C�c`t�4��+K�i�vr�?,ȷ-��� ��Q���1uo�M�iWͭ����F��k��\Zd=�	B0�x^�硣�~�D�*\��Fňh��v��$���d,ƌ��F�un<s6�C�>��o@w�9z��8��V'�@auJ�7B����2�
����@��q;�.EWFj!���H�@31��nȐ�y������΀���C��H1jH�XZ��V鳟�a��5>�m9�+x �_L�!�C�4_�nRbz�x��C��6�Q�����#�*���qTR~^"M#��kD�b��N'�=�����_7�T�&-xq`�D�i�z����'�/��((q�9�^�;n�6}�^��"b)t����+�e����Y�� ��$�9?mq=�$�u���F��X�ؗF.
�}s@j�t�pgH�$����y�.R"H�� M��F@?{����!q����J��@����ʷ�[�rQ :���$͍K���A�� �I�_��f��ԃ�"@S���C����δ�'˛�n�SD��:�@�	����4R3���q��8aϤ�p\�X'@u��{^�?K��7�� �i��]����AI���u� IHʗXD�?��\��s���ʭ�f��.ݏ��:����S0�3�ܥ��b%y�y��C
p�Ixxyvi���{�Rֶ��E��2²Ӱ��s�שh�b�6��[N�;�ي�m�w�R<3�[�fb;;N�o�Ou����(�D�@w��d�tNP�zWT�M4H +��K<��)�8@H)�F+Q?8��q�,^ס�q�
��(� c{;Ǉ�e�~w�[��`��0���s N"�S�a��lA�̷2���Xh����T�+QK`U��$�\����:`{�n	Lj��0X������<@ӈ���-�����~�$w�,�uq��3h�^���X+JB��=qD�1.��˗ᅵ�^n�.���؄�ו�o)���i�G?��O�EZ����+ w|��T��k������w��b���`�$��K��w�a3H�����1g�~��	�i[���n�<�D:=�������C�%n\/,/Z�e�̍�B���g���8c�o�z��>����
*�rj��;B�t��(`�Rg�1J�JX�g��]`�4�b<y�)�bB=dI�}�Gy���y�T����������5����G:Y��/��
"Ɔ� S�ca
"��b��*Os�e�^)�m���'��~4E��P�ۿ����De\�A8E��"bs�+p�W,��Ow��� �kj^�^�b9LS�U�����4ŏ32Ze�N`iY�L��5~� I!�(�� �1�J�BO�L�S��©�G1���xz��M���!b  �Sɋ�o�����wu�U�!��)�=Z<���8����β��s���+58�n
����F<��W�Jp�o���2n5��8��J{�{.�72�ZAWF~��ڗo�aq��)$4�G���d�h�	B���Gx��o���9�p�K�}f;}/d���{�f�Yw�����2�+�����n���~���Us��)����*H;6�!Pg���	h�{S��y�_�gn�l��+O|�z�@�R�$Ͼ�TZtz(�����tK��6=BT"�(H߂�3���bL��R�B=� S���,y!2�����e�+�mjA���*���ՕM	B�sv��6�o!��b���m>�.��<��+$��I�[����p���U]����K�0-i��gD�k�G<7b�40e��K߮6�_��b��v1�ؑ�v^�,�e�p�6O<<��SX�h
�9H�|H�eu�g#�[��^� L=�t����XhG#3��]H������!�y�7��ei����>�,���a����_�(�Vw̖J��,�4(��c�"�ӛ���xcnm!��L����k�s��o��|~�;Mdc&&�&j��0D̀�Hn=)��"#�6*o����<r��D$8���ڽIXr؇kgu3c��׷�2����� �&�CZwg����"X��^\z�F�4 `��O
gWy=ǘ�'I�W=�2ܛMDo��\�T| ��\��������R����n}�sQ�ιRMY
9ѐ���:aP��������y.�13���hG���6����TM���L�,��GJ���
^	�& U۴��7u����D�/���4�)D�,�F�>�%�D�N� �:����c&�j�Ѱ._�FZ��
��]�)���EX�%�D��Q�q).�3�ݍ�p�գ:#^�{Z��Xsɖ3���ac� � v���C~Ր����[c�����y�g&,)Ykئ�˅�>ճ���V{<s0Ӡ����5�r�)� 36�9f��1{VW
��5ܑ_#�J���`<��Xp�.>߄&��{�� �(e+�K:z�y�#dJ�� �@�/�mYb����/�}�8�a�H:y�rlQr��3dV�ڻr��6! ��a= ۬�K���}Vg�s�G�l�s����0����E�By�7��L=��Y,%����5GA���D�Hܮ$��M
��b@̚zYXHFVQɮQP]�/J�9Z$���\��4|Av���i����!b�M�J������v�HY������0���x��s�'8a�B���;�Ŋ�N+��"'O��i'�=a[��5!���4�jĭ�p����N�? ���B�����ѻdI̜�0YOl�Dhp!4|9�+i��P-R*���ߛ1e�Q��]C�R�P�'�p�.��k�4h]���J:0n�F�@vrF?ș�c�G �+����u�<OJY��T�:�%����6�k �P2��T�]��ܬ��G�w�(fᡛ�o���;a��ѼDT�Q�"3F~�У��pE��Ow�W��v#�{{O\k#�g�z{&R�C�|2�ͥ�OY5"j�߰�Kſ/�,�[f�:7+Z�_@��.�����/�_ x̋��^�TJ:MH�.U!��$��t�N�>6d(��<���v^�M�,�y����dbA��n� Gλ����ž��Sr��jM�#	bo0 ���ۢE[�6���<����%�i^���Ce��)�\��D��v`(W��e�Q�I�S�{��m��!h"�4�`,�����hѱ�9������ޙq�G8,w��"�N����x (ц�;�8U�VsX���7b���N���'��d��:i�Iq:���4�2���˥6�#m���;�t�\�	j�uRmU����g%�^(G������.��� �����ܔ0K��/K���Uг��:�M�#J��ዄPCzC�D_�2�m���zR ��%���
{X�۫{��l`'�V$o�Q�$�#P�-��0�i�YyL�y��Uf:
a�U:�Y6��YV�����[��^���8c�՞��C���G�d�EvJg�PƘ��� ��Ԅ��xV�<i�0(Kx�_�_⹸^]:bU�o�(d��>ߚ��괳q�F�8�PT��������<]#|��g%{�%��#�Kn�����8|G�HR�Y��ӏ��kbUT��'U�<��-
:[�l�\�ͷж[��6�X۹�"�t.C;�^�ުR:9���LY�^$(N��~��I��
�"	����"�a+�PMPG�y->f�Ql̜�xC����9!���i��I�B��������w2����M�����[�������P�ɀ�Fz�ER��9�łb��--nrLw������~�R�)kR�f�O��f�,�C�2s����������)�ERܮ;��{�vS�q�#�kG}hu����x���R]�AO-c�}��l�B��nSY�ZM+�������B�%5N�6>w|��~sr� pe�O��z�5C�}�II��؏V�>�J�	X�0	� $������VwٵV*F�C1��+�Cu�����&1. V�]���R�mLyF�:����Gj����6^�f+\�;v%��Y�����"q��%�/�����#G��ٮ��V�1zQk�c���1j��ndlzW�\��"� ��h2�BIr�s��[[Xܸ�'N��,c_C�.�c��j�kk����S���j���$�\�� 3���V���]��ee��+n�I��gnC�9�}��̅/Ά��U�m�1��l����`P^C�C���t\���]ҒR�PJ��E=�J�w�݃#���$
���f�Z���$H����]3t��?_T�-�rU.;�� �9Ǡ>2�|�BÒ���}1b���W���+o��>�V>R\��(S�[T�r�v�-}��Sm(rKn���+��I��TQ3�((�CL�6�����z��@ynD�z�0F*�t!���P�k��k����Qv"��b+������u��2"_c�:U}!��s�{����5��0��$Q�ZG��$�)��\��E����N�a1T#Ά_{�d��1�v��#�P��pih�����L�,�ǽ���FT���^%�(����b2�Z��4�N�����T6��!x�C��z/l���A�y���2��b�D/71�?Ƌ�X�����.De�'9�S*�9'�0t=���3o��^hK"I�����Ԛ ں�X>�2qs��pNO��ɫ�x�W�ͣ���7s߯1��T��a���� C�;?|�Kbঽ~��Ӻ�^z�'�i߾��!�O2P�d�X�8�Ȱ�m�ʗ�|��Ǆ�3�h|�Ic�}1���q����4jI��9Xk:�Ucp'��;�^<%��/cZ�w4����pqyL�+���VL5J�,u��_A)���ł?�G�2���R����aUw��ã�=��-�Y��h��9�iy��)�f�4)�'L�9��Mvp i�b�D6���E�Z�u�&�
��93���';�U*Q���:Enh����/yo����3�P�K�UC�j�(�P�L#)�m_�˕�R�:���j<�d�	�y���H��Kq��G��WBC��x$�7wty��T�X��o�Î0�݃)�;3{��V��ȫQ�P`e#�AeҾ	�����W"qC��h��R��-����i���#%�|S�F.�� 1�Կ�P� B7�DW��h��Kk{-�����ṃ�W~k��D��0��#P=�9��(~�I9����hn���� �}�咺�c%z�l�Zq�m_�n����H]*�����qL�(�0�=��Y�j��d��U�̓n�9%��T��mY��W����&.���c`����>��R�9"�I���=�It��S�	��\��R��g�e�?�;���4��u]tC�ɵL���
_�GMWRw<��������K=����eЄ�8d�"/�ɀ�-�l����y���E��T�h� �"8�e�?!��C(=����-�j��|��s�8l� �k7�[�>��}��V ��ՠ���\*{,��tI���-j-�.�S��1�d	7��^B/�<���C�1a.g�~������o��d(+ n��_5�95�H�� i	����T#��w�̌V����gײV�M���s񩧆�K���l["�1�u�&"��lH`1Sr�35
����9L|�.�cQ&����J��Š�*��g�#��!?��]q:���XM�;�mR�FX3��G��u��0{�N~�g�� $s,��������i��&��5�0���w�6luf��-�W8�`c��cA6��(Ga�����#˪�J����z[k ��PJ�s:��ޔQ�D��v�&�̾i�Z>JH������a�g�7&�}d�5k�N�z0ּA|,��+����5����S
��O�� �
����)n�-�(qyk�_�nG�İb�j �:����u8�T]�`�U�=����ĳM޵�ڵb���Ƴ�0Y���*�??z�6$"�jԼ���R��T]J�#\dX������MoZ���֘�z��G��pYuܚ��N4���Y��A�Ƈͯ��9Si4���._EQ[@���z��y��&�`7:/����י�,���q��T����-Vjq��K�}'E�V�ի���QZV?�$�%��J���9��!���{�xP���e�>e:��ů`~���(D~�-�������s�5��oܠ���1�2m�6�k�.,,
��j
��J~�#1�	W�b�F^��azi�K�,!�aL�<�����d����Ҿ�6���!XWx,	N�^A0'޹�_��wݵu��T7�0�B:i���� �^�'��J�=8�(�$�[bd'[tt����4��<��⚴��<�<+�\���_JO
"It �/���1z���M����F&�c���#�Տb8|z�ZZ8-0k)�yK�x5U��P�c�0?��,;ʰ��;�&�I_P�jS�w1��"������v�n��ܝ�A��:��}���4'��]�쭏$�'����M/玡t�Y�c�h�!��W˓(�V����@�A��co(Vݦ�$	��T^�^l�I{G�H�K����&"�5X���n,Qm!|�9����$�*ƭvG�nxF៟�_�]	p�H	���^�V����:n������p�NR�;������~MDi��|zt�7��U�	��V~#�{������NY� ��&���&8��y햻 ޿M�%�(Y�f2ɣ�9���.��w����q���)�J�U���H����}�y���Q���L�� V�t´�����%�E�e���S��.GoM@��Wn�=���N�A��o��g���(�,���u:�ECB���.m����#1?"�1t`<�/��s�a5�Y	ӎ�����׾���M�ȸnF�=�z鍉7����>QP��K2mI�(����@n�α���S�bv��ީ�0��h�f���i*0�s�	ko��7Q3��F��ap��ʹ݂�4�,򉯱��6�N�i�y�Kl�7���#�6*���ef�\LMq�
f�	$I��V�wL�@� �����z�e�ۃ��vm�� l
^�K��U���a0�b��k�X�,0�Ф���* :Ǚ�����/[9~���e^���vfYX��v��Q�'m�׸ԩ���j�����9�V!YM�F��� .��<#kz��t|��̄�"�g Q�M�jp8 '5�k�ɞ3	�z�ᒎ� �������4�)uĞ$G���	���~V��{���һ����;����Å��`�.)�u%��~4CT��8+�M�	)yas�pUe�;�-T�f�)G���&��S4��M^�;P�*j�B˕t_��e���f�tQA��'�B�v(���~�VA�YuyGиj��H�kA�G�Z��B�n*����c^,� �/���.c�c_��K�Ud�
 ���ZD}��d��=�h��E��X��*q�s�YhĭSːg����5d4�+�g�؍.'��vf?�{��"�v��k�ؖ%B���Xz/]ϗ�fxmj��U��7�O���H:��q� �`��݈LbjM}'�@�_�������@m��P	Vq�@�E�E*2��>�~	z������} vI�,�j�ߎ�Q�>F�h�24L�Wת��(�bq��9�z���
��	?焟����>�;��d��;��P�fمM��1b�)�w�ǥ��t!I���ޘ¦��UBg�g��t!�4�f�n����0(�O�>�?}�����1)%�D�ge�� u���JH��4�Uxf���o�O�j<{���_t
=X����Q5��;�<H@n���2ݳ�eGn������\��zz��N��yrߩ���<+Ҝ�8�v9,����b�b��d�1f6[�b>��Ď7�DL����q#�+�o�OQQ��`�{p��` 5�B}ϼ�0�,��u[ �щ���r�E�¸��q�"�0pf�!�����?�?��{�ye��s��k�ee��}��ס?��$]�x���_�~u\ة��Đ*E��w�6#���У=��F����\d�b��?����K,j����)�mL���HAp����c�-�jyeՆ���[�迍�����؞5jb��K��0��d��s�q������<��@� �QŒ
C7-��{�?�JW�w��2�!���B��˿w�w��Jc2|8��'�<`�D7��d���D��y2dpQ�iQe�MbR%�S5���,R�8��&���}\v�O#�'D(��]�_��E�])\[��e���%�o�*>< ??��T������f2]�����Y���_��Ԃz�<�"�D6'��/�â5z��K�*1�֗$���̗��w��y�.�y��?�l��9
4{.a�d4���׀j9�B ����+ �S?L�H�PF�;DM��Ȣ,���u��ӣKl��S,�OP��'���#�_��R�"7vܗ.'=�4��%r�1jM\�v��mZ����*�?GU��l3h���C>[�<�����د�䘋(��a�]�.��������s�	 �5y�^�����*��Z�A�J��s�k��_c�œM��h��`��x�&.7���Yeo��B3��A��݋ڇ��M�+��"S���zr�M@ʰ,M�c/=�X�a�	F��	.y�L)�� ��L��z��؅D/�bK'���f���O?=��7სǍ PY����O��RI���7j��_���v�v�9mS|�qRهO>�O>e]�c�Y��37m�~U̲���Ltg�$�Ý�By팪�� ���}���9�����Sf���$��*"����JՇ��� �ad6^-�;r�ӝh��請k�@��s����L�|~ĠC+D`��h�4����&vC�AOj��C�.�\����l"���Z����1�a�1�'�?Ó�b�G=�����l�sŘQ)F�)�����U�0�iС�Z@��O�?�QL/|LF��SX��6Nύ���*��^pۘ�Rll|���@�U(���*&���?�,�.�Qv�G�#�J�eR:z*����?��������U
�mM����A2�M���%�f�}~���:~�=)����^Rꠉ����a�'�OI�$r�^���a��݈�Թ4Lx�'x.fy�#ڂU���,0��0a���Ң�(��[��l3�m��k�g��3;U��4�\%7��f&��G�9�5u�J^�YWcS��sEn7�: ރ�5\�M��]Q���x�0� ��u	Q Ӣ;/�a㲧�
)#�-��C���<�4M`��u�J��� |�T� ^�)�� ���d[j���K}l�{W�4���R�Cw�A�"&��Y/�l��9Q_i�T 0�ig�C�M�2�B��5�I�V�ҭ������60fNw��2��OK���"o�)M�����M|⧣���6i�{*�G�i�]���r�fF@5�G8��cyQ�F����ĂY��=�!X� �� #�#��H5j�|y�s>�Y��%�1<凱xp�G�&��}�s���DKӓ{5R���P�jNT5���}�#���q�*���YVj��odA~����w��%����;A�2$k[����4�'�d��w� S�QH���D�I�6�lZLp�zPu��}&�_�����@����ڵ�f��K�3�}3F:;�U�y'�ޭ�t*-������5����Gn��]m���a�y�#Wv���d�<s�#gjǇ����?�[ _��_�:�2��*F��Q�d�z$�'����3��@����hcj5>$� ? ��H��f��ǸX��%�
z�@|>���UI�6�W\������7��S�=V#��4	��E�"�ªg:ӏm0Dv�ć��V?R�H
�,ʕ7u��e!�ؾ��'����8)��z5.6�^�.��t8��F>s���,У(�qG�x.��N��� ҩMA����|,�ښ�����-ae~�z��j-�&��ӯ�Bn�ӽ7r;�,�K��2h��Hw=��S�YϔrZv����Z��&x6x��O(��H�^x������/�$Pyp����6�b��ңo�F�[�cM;a�S-g�[�Y�'�Ϩ�S]v�1\ϡ���]�)��Ab�+߶YJ��lH ��Z��+���DY0e��=�!��&@T;2��*�¹nx��6H�R��p�ۣ\��Ĝ���-�IJ�dmԁ� 
�z ��$ׂTb!3
���!;��|{W�# m*v�p�@B�X`T�R7�wjX��fC1_Z��i9"�����Y#>�g����?�t\н:^'N��F��p}��R�h��O���)��ê4���M]+ܙ��i7�PS(��h�u������R�bwN�d=��c��%ϰ׍�3��˦*����?Qj��4�鸔"46��O�N� �\����_�O��+\�ul�q���H�l��*�¯u�q-�}�U ��"������.bxx�|��Pu�3M�Hԣ�be���������&�;�;qug���lgm}`~��.�@lR����,���>���P�\�qJ�g<u[�j^=��Ƽ��-C!�z#f�N=��W���V:�_�?���]j��ɶ���K���˵�s�	w��4aCS����l�������z��c}(c�m�:���B�%�kL��{��~�i�]�����f�N5��T�s܇�]v��}p��!��X#z���_����9�vn�u��hzêC{��yn�������{��&�1�RbCD<!}��x��N�d��$55t3G�4��3i"�������M����˴�W�'�Ъ�L�T|u���ȷ�^V BǇ���黔'*(sY��Mu�I�ǎ�?	.Ϲۼ:���>�M��~��U8�d��A�q�X�����a|�;�Y
�v"Z7,R��gwx�7 �W���
�2qe�h�V�%e4~�Hû���I�"�:{����ic�ǘ�����D<Y�F8��RL�"�ߐb�����)#6���˃�YDy
�7F���7|�C����d��6G��;B����2�\�{.�����8�b��? <g�Pͥ���+�h�<*R��_'F35-k��Xg����X����	�%v=dWWg�d�� vڲ�H^_��i��Ѝ����v앁%��}6���]	\��eK,��=)��5�S�A�#	�Y��[��P>bS�Q��9�j0r�qA�F����y��W�-�v	/۟������a��� >��q������@L�=*e�ع�7��T���.-�'S��P0.���ס�ےK��կθ�T��;��[��7���!������v���$j|Ѝf�����á�dӶ��$�!�������7��<�?��l1E��D�vJ��z���($�~ɳ%<���q�*e$��m��|�fk�}��J,���[]�ª}^Q���� �a�~vE�dm��}K.�>��PǙ+J�BNm>bS&,�l��#X�����'�����O =M�&��'ǳŌ��P�!��xV{�NU0��-�P��dϻ�iNI���zpޡ:g<ƿrk�I!�k�����ްf� �,W�F�N�?�8�`]�_�Ɗ�X�y|Y�Α^������Fl���4�q�����R��Q2BJi�D���	��yi4�e1�L��Y>{�Vŝ�:Q*��ܐ��uP}E��I��Uj�� H�̓�B��^"� 	~����(oX�ì����O�TlК��/��l�%1i�����ܦNH��%���2ky�XI�p�ܖ�3^�8D;��.6�c��2���mAq�*|���:?��2�I�~�I �"�x�#�� o�/�s��ȍ�+BI[Fw�L�w�U���L 0�N�.M�Yվ�57sh�a�!��<�
0�P=s�1�V-X�3_�.��#�ܙIϗ-���o���Y:Wl��$�N��h�}Z#�V��~�6�_\ �MSZ��-~G�Z�M��F�yF}	a������e+I�]5��)Jpֽ}͜�d*zQ쵟j������#��L�Qb�}3aKM�z�`���!t��|"5��o)�w��jz��9Q˚mZ�=zh->|]>,�5�����#C�"�{�8��s�?mʹ��xJ���U[K8��#2�U���).��w���+i�Q����u!喝ń�E��� K�L>t��p0��d�D���?���OL1�/ܩ|d<�ґ+� ��� Ԩ`s���̐?�d=�|4²��c�'5���(J!K;�hG��r�¾�:��2���TW���c�ڟSA�����m!j��H٨Qo�HK��gD"h/H��@Tp�ux�]�>ިwa���f%�hs��X�����/�|_=�Z�td��3��#�G�\`�ˏti�fD@���W�{d�Lj�ﺉ�}et��"�C�r�rH�U(����Ƥ^�N������a��ﶂ#K=��;6u��!�������ƌ��	t�?ew)����&�b�*��ʍPZu�>i9'�
�U�G���2����*}�q�T�D��H��y��ʷ��O`�K�SJ����O�����l�7J�5�x35���C]Ƴ=��@K���j?4x3�*`A�fq*s=�!�{�@a����Z��`�Ҕ�M�ܡ� >��x���(��aۍ��z�M��[����ƍ[%��B:�7cYE�87�M������(PXS&d���y�� ��U��.�#z���m;��W��~F7��:�Q8��[}��ɀ�窾��
�3����� �mLK8�a�/Ɯ� D�ˤ4�ܗ�����=+��7TM�K��r;G_L���T�xqɼ�`��HI�w�u�7�7��["s,��_�>3�~����,E�E��7th���!G0�~pt�iD?ծK$bg�g�r�{DMΝs2�Y/�W��A��c�x�Z�ጬ�`�[}-��[�8�=e�R��8�99�EN҉詈!N����`	d/ɰ�<ÚpV=�j9֜e(�u�?��/7-�s�":����_ k��$D@ ��ʡq�=Y؅�pcd�Ovb'���&͛՟�� ����9t�eu��g�$� ������LU�S�j�[С���Zos������@�pF{fu,�SC�U�C�W0����'�޲�����JvM@B"E5�� �W�� �Ԕ�l���6��;��ia}�5�>�E���Cf-p�������lh?%v�M�lO��l�4_z�Ϡ� د�NNҾ�X��TV*-U6u�S�������K����+�L����PuE��M�t���Ha�������x�@�&="���yKC\2�v:��w��7\��g�C���#+��`&�ܙƁ������a5*.����m� Xsm��������'��S�bC?xb��o{��YEḴ��v�e���p�e[��©��_���u�6'�e�=nFnv��e����Nc �E���!XU$}��"���\H�5y_%-xٜ��^��H�=�ϝ2v&�!�@���s��3hh $c
�y_[!,b�֯8�"U�ovɛ�a2�������{�&F�Q����Jx;���&��=�T|��h��j=�E,����R����WԳ��&Yɠ"������Љ��_�����S��y��D̍�mO1���bN�QS�����?SZt����`׊������#��D�	x��L��fU9�G�I%ĽS�3ύCq�{:�o�����bϦ�����=�a؈��X�}��2�Ɍ�
L	b�!��\�|���c�y�e��{��`�t��^�Ec��
�~�i0U�#�gy!�ʐ�x���Xd>�Yr���,J��������)���ŉ+d��������|�L�/�b*��\4�S�����DnL�]k,��пד����j\��U�ES2M���;S���f*��z9ׂH+�<�&�$�f�i��me���&��slv����3��
tzty"����EK!��D�f8�ҳhpc/v�Y �s��_�:�H�Q��?�+��(�)64����՜8��2�;
���-|��*��#���GU����T8#}����kC�l�^���ob9��Ζ�e�|9�]����&�hIpf�)��elbz3�)#0]�W&���
r��{��T���%�u2e��W=R�񻗜6A�XcpC1BI�@
ŉ�K����Z/	y�W�� ����.��m[iw7�1���]�"�4��r����
���Y��^�:K2���L{�%�ao��9��@,3���c���Qv�,��k�N���-��ު8��9���˶�TϽXU`�:��	W��H)�b���T�}�m:q\s�]@#����N�lR�LȂ���ds#}���*���>~��� ��d,���P=��2�3ܫ��9R!HJn�6R���I�IQ�˧��	��V�7F4M�?m���\�FE��V�<~��/	W7��Uc7���ӊ�%u��8h9ǃT#�b�هbb[K�S�{�=�<,��d��	����I�"� $N0o�{z�ȕz���'f���S�w�C����/��4�]usL���¹6�S�xe�W�Ȩ�e^��lXG�2�˺ѦC[p\R�@�La�⩵us�����Tζ���Cޮ�c>��za��Bf�8��^q�:Ĩ
V��w�����y���* �vclQ����5�4�z�u�7���Joʽ�J�W���������t�u����p�����G��c���z԰:��M��M%��h����!c��'�����L�s�3��-�w�qL��c��Y���V��mf2a^`��RO©�B��gA�-�7<�ѻ��o�م��}�QU\U�8f���{�BZ�]� {���^g����Yk6Ͼ6�7�߷+"C����Īp����