
module DE2_115_SOPC (
	clk_clk,
	reset_reset_n,
	pio_led_external_connection_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[7:0]	pio_led_external_connection_export;
endmodule
