-- megafunction wizard: %LPM_ADD_SUB%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: lpm_add_sub 

-- ============================================================
-- File Name: wb_audioStream_channelAdder.vhd
-- Megafunction Name(s):
-- 			lpm_add_sub
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 8.0 Build 231 07/10/2008 SP 1 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2008 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY lpm;
USE lpm.all;

ENTITY wb_audioStream_channelAdder IS
	PORT
	(
		dataa		: IN STD_LOGIC_VECTOR (16 DOWNTO 0);
		datab		: IN STD_LOGIC_VECTOR (16 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (16 DOWNTO 0)
	);
END wb_audioStream_channelAdder;


ARCHITECTURE SYN OF wb_audiostream_channeladder IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (16 DOWNTO 0);



	COMPONENT lpm_add_sub
	GENERIC (
		lpm_direction		: STRING;
		lpm_hint		: STRING;
		lpm_representation		: STRING;
		lpm_type		: STRING;
		lpm_width		: NATURAL
	);
	PORT (
			dataa	: IN STD_LOGIC_VECTOR (16 DOWNTO 0);
			datab	: IN STD_LOGIC_VECTOR (16 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (16 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(16 DOWNTO 0);

	lpm_add_sub_component : lpm_add_sub
	GENERIC MAP (
		lpm_direction => "ADD",
		lpm_hint => "ONE_INPUT_IS_CONSTANT=NO,CIN_USED=NO,CBX_MODULE_PREFIX=wb_audioStream_channelAdder",
		lpm_representation => "SIGNED",
		lpm_type => "LPM_ADD_SUB",
		lpm_width => 17
	)
	PORT MAP (
		dataa => dataa,
		datab => datab,
		result => sub_wire0
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: CarryIn NUMERIC "0"
-- Retrieval info: PRIVATE: CarryOut NUMERIC "0"
-- Retrieval info: PRIVATE: ConstantA NUMERIC "0"
-- Retrieval info: PRIVATE: ConstantB NUMERIC "0"
-- Retrieval info: PRIVATE: Function NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
-- Retrieval info: PRIVATE: LPM_PIPELINE NUMERIC "0"
-- Retrieval info: PRIVATE: Latency NUMERIC "0"
-- Retrieval info: PRIVATE: Overflow NUMERIC "0"
-- Retrieval info: PRIVATE: RadixA NUMERIC "10"
-- Retrieval info: PRIVATE: RadixB NUMERIC "10"
-- Retrieval info: PRIVATE: Representation NUMERIC "0"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: ValidCtA NUMERIC "0"
-- Retrieval info: PRIVATE: ValidCtB NUMERIC "0"
-- Retrieval info: PRIVATE: WhichConstant NUMERIC "0"
-- Retrieval info: PRIVATE: aclr NUMERIC "0"
-- Retrieval info: PRIVATE: clken NUMERIC "0"
-- Retrieval info: PRIVATE: nBit NUMERIC "17"
-- Retrieval info: CONSTANT: LPM_DIRECTION STRING "ADD"
-- Retrieval info: CONSTANT: LPM_HINT STRING "ONE_INPUT_IS_CONSTANT=NO,CIN_USED=NO"
-- Retrieval info: CONSTANT: LPM_REPRESENTATION STRING "SIGNED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_ADD_SUB"
-- Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "17"
-- Retrieval info: USED_PORT: dataa 0 0 17 0 INPUT NODEFVAL dataa[16..0]
-- Retrieval info: USED_PORT: datab 0 0 17 0 INPUT NODEFVAL datab[16..0]
-- Retrieval info: USED_PORT: result 0 0 17 0 OUTPUT NODEFVAL result[16..0]
-- Retrieval info: CONNECT: result 0 0 17 0 @result 0 0 17 0
-- Retrieval info: CONNECT: @dataa 0 0 17 0 dataa 0 0 17 0
-- Retrieval info: CONNECT: @datab 0 0 17 0 datab 0 0 17 0
-- Retrieval info: LIBRARY: lpm lpm.lpm_components.all
-- Retrieval info: GEN_FILE: TYPE_NORMAL wb_audioStream_channelAdder.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL wb_audioStream_channelAdder.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL wb_audioStream_channelAdder.cmp FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL wb_audioStream_channelAdder.bsf TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL wb_audioStream_channelAdder_inst.vhd FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL wb_audioStream_channelAdder_waveforms.html FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL wb_audioStream_channelAdder_wave*.jpg FALSE
-- Retrieval info: LIB_FILE: lpm
-- Retrieval info: CBX_MODULE_PREFIX: ON
